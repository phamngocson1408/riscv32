module MulAddRecFNToRaw_postMul( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190483.2]
  input         io_fromPreMul_isSigNaNAny, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_isNaNAOrB, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_isInfA, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_isZeroA, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_isInfB, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_isZeroB, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_signProd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_isNaNC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_isInfC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_isZeroC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input  [9:0]  io_fromPreMul_sExpSum, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_doSubMags, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_CIsDominant, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input  [4:0]  io_fromPreMul_CDom_CAlignDist, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input  [25:0] io_fromPreMul_highAlignedSigC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input         io_fromPreMul_bit0AlignedSigC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input  [48:0] io_mulAddResult, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  input  [2:0]  io_roundingMode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  output        io_invalidExc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  output        io_rawOut_isNaN, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  output        io_rawOut_isInf, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  output        io_rawOut_isZero, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  output        io_rawOut_sign, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  output [9:0]  io_rawOut_sExp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
  output [26:0] io_rawOut_sig // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190484.4]
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45:freechips.rocketchip.system.DefaultRV32Config.fir@190487.4]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42:freechips.rocketchip.system.DefaultRV32Config.fir@190488.4]
  wire [25:0] _T_2; // @[MulAddRecFN.scala 195:47:freechips.rocketchip.system.DefaultRV32Config.fir@190491.4]
  wire [25:0] _T_3; // @[MulAddRecFN.scala 194:16:freechips.rocketchip.system.DefaultRV32Config.fir@190492.4]
  wire [74:0] sigSum; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190495.4]
  wire [1:0] _T_6; // @[MulAddRecFN.scala 205:69:freechips.rocketchip.system.DefaultRV32Config.fir@190496.4]
  wire [9:0] _GEN_0; // @[MulAddRecFN.scala 205:43:freechips.rocketchip.system.DefaultRV32Config.fir@190497.4]
  wire [9:0] CDom_sExp; // @[MulAddRecFN.scala 205:43:freechips.rocketchip.system.DefaultRV32Config.fir@190499.4]
  wire [49:0] _T_10; // @[MulAddRecFN.scala 208:13:freechips.rocketchip.system.DefaultRV32Config.fir@190501.4]
  wire [49:0] _T_14; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190505.4]
  wire [49:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12:freechips.rocketchip.system.DefaultRV32Config.fir@190506.4]
  wire [23:0] _T_16; // @[MulAddRecFN.scala 217:14:freechips.rocketchip.system.DefaultRV32Config.fir@190508.4]
  wire  _T_17; // @[MulAddRecFN.scala 217:36:freechips.rocketchip.system.DefaultRV32Config.fir@190509.4]
  wire  _T_19; // @[MulAddRecFN.scala 218:37:freechips.rocketchip.system.DefaultRV32Config.fir@190511.4]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12:freechips.rocketchip.system.DefaultRV32Config.fir@190512.4]
  wire [80:0] _GEN_1; // @[MulAddRecFN.scala 221:24:freechips.rocketchip.system.DefaultRV32Config.fir@190513.4]
  wire [80:0] _T_20; // @[MulAddRecFN.scala 221:24:freechips.rocketchip.system.DefaultRV32Config.fir@190513.4]
  wire [28:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56:freechips.rocketchip.system.DefaultRV32Config.fir@190514.4]
  wire [26:0] in_orReduceBy4; // @[MulAddRecFN.scala 224:53:freechips.rocketchip.system.DefaultRV32Config.fir@190516.4]
  wire  reducedVec_orReduceBy4_0; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190520.4]
  wire  reducedVec_orReduceBy4_1; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190523.4]
  wire  reducedVec_orReduceBy4_2; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190526.4]
  wire  reducedVec_orReduceBy4_3; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190529.4]
  wire  reducedVec_orReduceBy4_4; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190532.4]
  wire  reducedVec_orReduceBy4_5; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190535.4]
  wire  reducedVec_orReduceBy4_6; // @[primitives.scala 212:57:freechips.rocketchip.system.DefaultRV32Config.fir@190538.4]
  wire [6:0] _T_41; // @[primitives.scala 213:20:freechips.rocketchip.system.DefaultRV32Config.fir@190545.4]
  wire [2:0] in_inv; // @[primitives.scala 118:30:freechips.rocketchip.system.DefaultRV32Config.fir@190547.4]
  wire [8:0] shift; // @[primitives.scala 160:58:freechips.rocketchip.system.DefaultRV32Config.fir@190548.4]
  wire [5:0] my_lowMask_1; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190564.4]
  wire [6:0] _GEN_2; // @[MulAddRecFN.scala 224:72:freechips.rocketchip.system.DefaultRV32Config.fir@190565.4]
  wire [6:0] _T_58; // @[MulAddRecFN.scala 224:72:freechips.rocketchip.system.DefaultRV32Config.fir@190565.4]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73:freechips.rocketchip.system.DefaultRV32Config.fir@190566.4]
  wire  _T_61; // @[MulAddRecFN.scala 228:32:freechips.rocketchip.system.DefaultRV32Config.fir@190569.4]
  wire  _T_62; // @[MulAddRecFN.scala 228:36:freechips.rocketchip.system.DefaultRV32Config.fir@190570.4]
  wire  _T_63; // @[MulAddRecFN.scala 228:61:freechips.rocketchip.system.DefaultRV32Config.fir@190571.4]
  wire [26:0] CDom_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190572.4]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36:freechips.rocketchip.system.DefaultRV32Config.fir@190573.4]
  wire [50:0] _T_65; // @[MulAddRecFN.scala 237:13:freechips.rocketchip.system.DefaultRV32Config.fir@190575.4]
  wire [50:0] _GEN_3; // @[MulAddRecFN.scala 238:41:freechips.rocketchip.system.DefaultRV32Config.fir@190577.4]
  wire [50:0] _T_68; // @[MulAddRecFN.scala 238:41:freechips.rocketchip.system.DefaultRV32Config.fir@190578.4]
  wire [50:0] in_orReduceBy2; // @[MulAddRecFN.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@190579.4]
  wire  reducedVec_orReduceBy2__0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190583.4]
  wire  reducedVec_orReduceBy2__1; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190586.4]
  wire  reducedVec_orReduceBy2__2; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190589.4]
  wire  reducedVec_orReduceBy2__3; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190592.4]
  wire  reducedVec_orReduceBy2__4; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190595.4]
  wire  reducedVec_orReduceBy2__5; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190598.4]
  wire  reducedVec_orReduceBy2__6; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190601.4]
  wire  reducedVec_orReduceBy2__7; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190604.4]
  wire  reducedVec_orReduceBy2__8; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190607.4]
  wire  reducedVec_orReduceBy2__9; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190610.4]
  wire  reducedVec_orReduceBy2__10; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190613.4]
  wire  reducedVec_orReduceBy2__11; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190616.4]
  wire  reducedVec_orReduceBy2__12; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190619.4]
  wire  reducedVec_orReduceBy2__13; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190622.4]
  wire  reducedVec_orReduceBy2__14; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190625.4]
  wire  reducedVec_orReduceBy2__15; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190628.4]
  wire  reducedVec_orReduceBy2__16; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190631.4]
  wire  reducedVec_orReduceBy2__17; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190634.4]
  wire  reducedVec_orReduceBy2__18; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190637.4]
  wire  reducedVec_orReduceBy2__19; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190640.4]
  wire  reducedVec_orReduceBy2__20; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190643.4]
  wire  reducedVec_orReduceBy2__21; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190646.4]
  wire  reducedVec_orReduceBy2__22; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190649.4]
  wire  reducedVec_orReduceBy2__23; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190652.4]
  wire  reducedVec_orReduceBy2__24; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190655.4]
  wire  reducedVec_orReduceBy2__25; // @[primitives.scala 193:15:freechips.rocketchip.system.DefaultRV32Config.fir@190657.4]
  wire [5:0] _T_125; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190664.4]
  wire [12:0] _T_132; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190671.4]
  wire [5:0] _T_137; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190676.4]
  wire [25:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190684.4]
  wire [4:0] _T_171; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190711.4]
  wire [4:0] _T_172; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190712.4]
  wire [4:0] _T_173; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190713.4]
  wire [4:0] _T_174; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190714.4]
  wire [4:0] _T_175; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190715.4]
  wire [4:0] _T_176; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190716.4]
  wire [4:0] _T_177; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190717.4]
  wire [4:0] _T_178; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190718.4]
  wire [4:0] _T_179; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190719.4]
  wire [4:0] _T_180; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190720.4]
  wire [4:0] _T_181; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190721.4]
  wire [4:0] _T_182; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190722.4]
  wire [4:0] _T_183; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190723.4]
  wire [4:0] _T_184; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190724.4]
  wire [4:0] _T_185; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190725.4]
  wire [4:0] _T_186; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190726.4]
  wire [4:0] _T_187; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190727.4]
  wire [4:0] _T_188; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190728.4]
  wire [4:0] _T_189; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190729.4]
  wire [4:0] _T_190; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190730.4]
  wire [4:0] _T_191; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190731.4]
  wire [4:0] _T_192; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190732.4]
  wire [4:0] _T_193; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190733.4]
  wire [4:0] _T_194; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190734.4]
  wire [4:0] notCDom_normDistReduced2; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190735.4]
  wire [5:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56:freechips.rocketchip.system.DefaultRV32Config.fir@190736.4]
  wire [6:0] _T_195; // @[MulAddRecFN.scala 243:69:freechips.rocketchip.system.DefaultRV32Config.fir@190737.4]
  wire [9:0] _GEN_4; // @[MulAddRecFN.scala 243:46:freechips.rocketchip.system.DefaultRV32Config.fir@190738.4]
  wire [9:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46:freechips.rocketchip.system.DefaultRV32Config.fir@190740.4]
  wire [113:0] _GEN_5; // @[MulAddRecFN.scala 245:27:freechips.rocketchip.system.DefaultRV32Config.fir@190741.4]
  wire [113:0] _T_198; // @[MulAddRecFN.scala 245:27:freechips.rocketchip.system.DefaultRV32Config.fir@190741.4]
  wire [28:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50:freechips.rocketchip.system.DefaultRV32Config.fir@190742.4]
  wire [12:0] in_orReduceBy2_1; // @[MulAddRecFN.scala 249:39:freechips.rocketchip.system.DefaultRV32Config.fir@190743.4]
  wire  reducedVec_orReduceBy2_1_0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190748.4]
  wire  reducedVec_orReduceBy2_1_1; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190751.4]
  wire  reducedVec_orReduceBy2_1_2; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190754.4]
  wire  reducedVec_orReduceBy2_1_3; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190757.4]
  wire  reducedVec_orReduceBy2_1_4; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190760.4]
  wire  reducedVec_orReduceBy2_1_5; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190763.4]
  wire  reducedVec_orReduceBy2_1_6; // @[primitives.scala 193:15:freechips.rocketchip.system.DefaultRV32Config.fir@190765.4]
  wire [6:0] _T_219; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190773.4]
  wire [3:0] in_inv_1; // @[primitives.scala 118:30:freechips.rocketchip.system.DefaultRV32Config.fir@190775.4]
  wire [16:0] shift_1; // @[primitives.scala 160:58:freechips.rocketchip.system.DefaultRV32Config.fir@190776.4]
  wire [5:0] my_lowMask_1_1; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190792.4]
  wire [6:0] _GEN_6; // @[MulAddRecFN.scala 249:78:freechips.rocketchip.system.DefaultRV32Config.fir@190793.4]
  wire [6:0] _T_236; // @[MulAddRecFN.scala 249:78:freechips.rocketchip.system.DefaultRV32Config.fir@190793.4]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11:freechips.rocketchip.system.DefaultRV32Config.fir@190794.4]
  wire  _T_239; // @[MulAddRecFN.scala 254:35:freechips.rocketchip.system.DefaultRV32Config.fir@190797.4]
  wire  _T_240; // @[MulAddRecFN.scala 254:39:freechips.rocketchip.system.DefaultRV32Config.fir@190798.4]
  wire [26:0] notCDom_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190799.4]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50:freechips.rocketchip.system.DefaultRV32Config.fir@190801.4]
  wire  _T_242; // @[MulAddRecFN.scala 261:36:freechips.rocketchip.system.DefaultRV32Config.fir@190802.4]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12:freechips.rocketchip.system.DefaultRV32Config.fir@190803.4]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49:freechips.rocketchip.system.DefaultRV32Config.fir@190804.4]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44:freechips.rocketchip.system.DefaultRV32Config.fir@190805.4]
  wire  _T_243; // @[MulAddRecFN.scala 269:32:freechips.rocketchip.system.DefaultRV32Config.fir@190806.4]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58:freechips.rocketchip.system.DefaultRV32Config.fir@190807.4]
  wire  _T_244; // @[MulAddRecFN.scala 274:31:freechips.rocketchip.system.DefaultRV32Config.fir@190808.4]
  wire  _T_245; // @[MulAddRecFN.scala 273:35:freechips.rocketchip.system.DefaultRV32Config.fir@190809.4]
  wire  _T_246; // @[MulAddRecFN.scala 275:32:freechips.rocketchip.system.DefaultRV32Config.fir@190810.4]
  wire  _T_247; // @[MulAddRecFN.scala 274:57:freechips.rocketchip.system.DefaultRV32Config.fir@190811.4]
  wire  _T_248; // @[MulAddRecFN.scala 276:10:freechips.rocketchip.system.DefaultRV32Config.fir@190812.4]
  wire  _T_250; // @[MulAddRecFN.scala 276:36:freechips.rocketchip.system.DefaultRV32Config.fir@190814.4]
  wire  _T_251; // @[MulAddRecFN.scala 277:61:freechips.rocketchip.system.DefaultRV32Config.fir@190815.4]
  wire  _T_252; // @[MulAddRecFN.scala 278:35:freechips.rocketchip.system.DefaultRV32Config.fir@190816.4]
  wire  _T_255; // @[MulAddRecFN.scala 285:14:freechips.rocketchip.system.DefaultRV32Config.fir@190822.4]
  wire  _T_256; // @[MulAddRecFN.scala 285:42:freechips.rocketchip.system.DefaultRV32Config.fir@190823.4]
  wire  _T_258; // @[MulAddRecFN.scala 287:27:freechips.rocketchip.system.DefaultRV32Config.fir@190826.4]
  wire  _T_259; // @[MulAddRecFN.scala 288:31:freechips.rocketchip.system.DefaultRV32Config.fir@190827.4]
  wire  _T_260; // @[MulAddRecFN.scala 287:54:freechips.rocketchip.system.DefaultRV32Config.fir@190828.4]
  wire  _T_261; // @[MulAddRecFN.scala 289:29:freechips.rocketchip.system.DefaultRV32Config.fir@190829.4]
  wire  _T_262; // @[MulAddRecFN.scala 289:26:freechips.rocketchip.system.DefaultRV32Config.fir@190830.4]
  wire  _T_263; // @[MulAddRecFN.scala 289:48:freechips.rocketchip.system.DefaultRV32Config.fir@190831.4]
  wire  _T_264; // @[MulAddRecFN.scala 290:36:freechips.rocketchip.system.DefaultRV32Config.fir@190832.4]
  wire  _T_265; // @[MulAddRecFN.scala 288:43:freechips.rocketchip.system.DefaultRV32Config.fir@190833.4]
  wire  _T_266; // @[MulAddRecFN.scala 291:26:freechips.rocketchip.system.DefaultRV32Config.fir@190834.4]
  wire  _T_267; // @[MulAddRecFN.scala 292:37:freechips.rocketchip.system.DefaultRV32Config.fir@190835.4]
  wire  _T_268; // @[MulAddRecFN.scala 291:46:freechips.rocketchip.system.DefaultRV32Config.fir@190836.4]
  wire  _T_269; // @[MulAddRecFN.scala 290:48:freechips.rocketchip.system.DefaultRV32Config.fir@190837.4]
  wire  _T_270; // @[MulAddRecFN.scala 293:10:freechips.rocketchip.system.DefaultRV32Config.fir@190838.4]
  wire  _T_271; // @[MulAddRecFN.scala 293:31:freechips.rocketchip.system.DefaultRV32Config.fir@190839.4]
  wire  _T_272; // @[MulAddRecFN.scala 293:28:freechips.rocketchip.system.DefaultRV32Config.fir@190840.4]
  wire  _T_273; // @[MulAddRecFN.scala 294:17:freechips.rocketchip.system.DefaultRV32Config.fir@190841.4]
  wire  _T_274; // @[MulAddRecFN.scala 293:49:freechips.rocketchip.system.DefaultRV32Config.fir@190842.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45:freechips.rocketchip.system.DefaultRV32Config.fir@190487.4]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42:freechips.rocketchip.system.DefaultRV32Config.fir@190488.4]
  assign _T_2 = io_fromPreMul_highAlignedSigC + 26'h1; // @[MulAddRecFN.scala 195:47:freechips.rocketchip.system.DefaultRV32Config.fir@190491.4]
  assign _T_3 = io_mulAddResult[48] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16:freechips.rocketchip.system.DefaultRV32Config.fir@190492.4]
  assign sigSum = {_T_3,io_mulAddResult[47:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190495.4]
  assign _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69:freechips.rocketchip.system.DefaultRV32Config.fir@190496.4]
  assign _GEN_0 = {{8{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43:freechips.rocketchip.system.DefaultRV32Config.fir@190497.4]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43:freechips.rocketchip.system.DefaultRV32Config.fir@190499.4]
  assign _T_10 = ~sigSum[74:25]; // @[MulAddRecFN.scala 208:13:freechips.rocketchip.system.DefaultRV32Config.fir@190501.4]
  assign _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[25:24],sigSum[72:26]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190505.4]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? _T_10 : _T_14; // @[MulAddRecFN.scala 207:12:freechips.rocketchip.system.DefaultRV32Config.fir@190506.4]
  assign _T_16 = ~sigSum[24:1]; // @[MulAddRecFN.scala 217:14:freechips.rocketchip.system.DefaultRV32Config.fir@190508.4]
  assign _T_17 = _T_16 != 24'h0; // @[MulAddRecFN.scala 217:36:freechips.rocketchip.system.DefaultRV32Config.fir@190509.4]
  assign _T_19 = sigSum[25:1] != 25'h0; // @[MulAddRecFN.scala 218:37:freechips.rocketchip.system.DefaultRV32Config.fir@190511.4]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12:freechips.rocketchip.system.DefaultRV32Config.fir@190512.4]
  assign _GEN_1 = {{31'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24:freechips.rocketchip.system.DefaultRV32Config.fir@190513.4]
  assign _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24:freechips.rocketchip.system.DefaultRV32Config.fir@190513.4]
  assign CDom_mainSig = _T_20[49:21]; // @[MulAddRecFN.scala 221:56:freechips.rocketchip.system.DefaultRV32Config.fir@190514.4]
  assign in_orReduceBy4 = {CDom_absSigSum[23:0], 3'h0}; // @[MulAddRecFN.scala 224:53:freechips.rocketchip.system.DefaultRV32Config.fir@190516.4]
  assign reducedVec_orReduceBy4_0 = in_orReduceBy4[3:0] != 4'h0; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190520.4]
  assign reducedVec_orReduceBy4_1 = in_orReduceBy4[7:4] != 4'h0; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190523.4]
  assign reducedVec_orReduceBy4_2 = in_orReduceBy4[11:8] != 4'h0; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190526.4]
  assign reducedVec_orReduceBy4_3 = in_orReduceBy4[15:12] != 4'h0; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190529.4]
  assign reducedVec_orReduceBy4_4 = in_orReduceBy4[19:16] != 4'h0; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190532.4]
  assign reducedVec_orReduceBy4_5 = in_orReduceBy4[23:20] != 4'h0; // @[primitives.scala 209:54:freechips.rocketchip.system.DefaultRV32Config.fir@190535.4]
  assign reducedVec_orReduceBy4_6 = in_orReduceBy4[26:24] != 3'h0; // @[primitives.scala 212:57:freechips.rocketchip.system.DefaultRV32Config.fir@190538.4]
  assign _T_41 = {reducedVec_orReduceBy4_6,reducedVec_orReduceBy4_5,reducedVec_orReduceBy4_4,reducedVec_orReduceBy4_3,reducedVec_orReduceBy4_2,reducedVec_orReduceBy4_1,reducedVec_orReduceBy4_0}; // @[primitives.scala 213:20:freechips.rocketchip.system.DefaultRV32Config.fir@190545.4]
  assign in_inv = ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[primitives.scala 118:30:freechips.rocketchip.system.DefaultRV32Config.fir@190547.4]
  assign shift = -9'sh100 >>> in_inv; // @[primitives.scala 160:58:freechips.rocketchip.system.DefaultRV32Config.fir@190548.4]
  assign my_lowMask_1 = {shift[1],shift[2],shift[3],shift[4],shift[5],shift[6]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190564.4]
  assign _GEN_2 = {{1'd0}, my_lowMask_1}; // @[MulAddRecFN.scala 224:72:freechips.rocketchip.system.DefaultRV32Config.fir@190565.4]
  assign _T_58 = _T_41 & _GEN_2; // @[MulAddRecFN.scala 224:72:freechips.rocketchip.system.DefaultRV32Config.fir@190565.4]
  assign CDom_reduced4SigExtra = _T_58 != 7'h0; // @[MulAddRecFN.scala 225:73:freechips.rocketchip.system.DefaultRV32Config.fir@190566.4]
  assign _T_61 = CDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 228:32:freechips.rocketchip.system.DefaultRV32Config.fir@190569.4]
  assign _T_62 = _T_61 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36:freechips.rocketchip.system.DefaultRV32Config.fir@190570.4]
  assign _T_63 = _T_62 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61:freechips.rocketchip.system.DefaultRV32Config.fir@190571.4]
  assign CDom_sig = {CDom_mainSig[28:3],_T_63}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190572.4]
  assign notCDom_signSigSum = sigSum[51]; // @[MulAddRecFN.scala 234:36:freechips.rocketchip.system.DefaultRV32Config.fir@190573.4]
  assign _T_65 = ~sigSum[50:0]; // @[MulAddRecFN.scala 237:13:freechips.rocketchip.system.DefaultRV32Config.fir@190575.4]
  assign _GEN_3 = {{50'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41:freechips.rocketchip.system.DefaultRV32Config.fir@190577.4]
  assign _T_68 = sigSum[50:0] + _GEN_3; // @[MulAddRecFN.scala 238:41:freechips.rocketchip.system.DefaultRV32Config.fir@190578.4]
  assign in_orReduceBy2 = notCDom_signSigSum ? _T_65 : _T_68; // @[MulAddRecFN.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@190579.4]
  assign reducedVec_orReduceBy2__0 = in_orReduceBy2[1:0] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190583.4]
  assign reducedVec_orReduceBy2__1 = in_orReduceBy2[3:2] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190586.4]
  assign reducedVec_orReduceBy2__2 = in_orReduceBy2[5:4] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190589.4]
  assign reducedVec_orReduceBy2__3 = in_orReduceBy2[7:6] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190592.4]
  assign reducedVec_orReduceBy2__4 = in_orReduceBy2[9:8] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190595.4]
  assign reducedVec_orReduceBy2__5 = in_orReduceBy2[11:10] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190598.4]
  assign reducedVec_orReduceBy2__6 = in_orReduceBy2[13:12] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190601.4]
  assign reducedVec_orReduceBy2__7 = in_orReduceBy2[15:14] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190604.4]
  assign reducedVec_orReduceBy2__8 = in_orReduceBy2[17:16] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190607.4]
  assign reducedVec_orReduceBy2__9 = in_orReduceBy2[19:18] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190610.4]
  assign reducedVec_orReduceBy2__10 = in_orReduceBy2[21:20] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190613.4]
  assign reducedVec_orReduceBy2__11 = in_orReduceBy2[23:22] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190616.4]
  assign reducedVec_orReduceBy2__12 = in_orReduceBy2[25:24] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190619.4]
  assign reducedVec_orReduceBy2__13 = in_orReduceBy2[27:26] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190622.4]
  assign reducedVec_orReduceBy2__14 = in_orReduceBy2[29:28] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190625.4]
  assign reducedVec_orReduceBy2__15 = in_orReduceBy2[31:30] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190628.4]
  assign reducedVec_orReduceBy2__16 = in_orReduceBy2[33:32] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190631.4]
  assign reducedVec_orReduceBy2__17 = in_orReduceBy2[35:34] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190634.4]
  assign reducedVec_orReduceBy2__18 = in_orReduceBy2[37:36] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190637.4]
  assign reducedVec_orReduceBy2__19 = in_orReduceBy2[39:38] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190640.4]
  assign reducedVec_orReduceBy2__20 = in_orReduceBy2[41:40] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190643.4]
  assign reducedVec_orReduceBy2__21 = in_orReduceBy2[43:42] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190646.4]
  assign reducedVec_orReduceBy2__22 = in_orReduceBy2[45:44] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190649.4]
  assign reducedVec_orReduceBy2__23 = in_orReduceBy2[47:46] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190652.4]
  assign reducedVec_orReduceBy2__24 = in_orReduceBy2[49:48] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190655.4]
  assign reducedVec_orReduceBy2__25 = in_orReduceBy2[50]; // @[primitives.scala 193:15:freechips.rocketchip.system.DefaultRV32Config.fir@190657.4]
  assign _T_125 = {reducedVec_orReduceBy2__5,reducedVec_orReduceBy2__4,reducedVec_orReduceBy2__3,reducedVec_orReduceBy2__2,reducedVec_orReduceBy2__1,reducedVec_orReduceBy2__0}; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190664.4]
  assign _T_132 = {reducedVec_orReduceBy2__12,reducedVec_orReduceBy2__11,reducedVec_orReduceBy2__10,reducedVec_orReduceBy2__9,reducedVec_orReduceBy2__8,reducedVec_orReduceBy2__7,reducedVec_orReduceBy2__6,_T_125}; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190671.4]
  assign _T_137 = {reducedVec_orReduceBy2__18,reducedVec_orReduceBy2__17,reducedVec_orReduceBy2__16,reducedVec_orReduceBy2__15,reducedVec_orReduceBy2__14,reducedVec_orReduceBy2__13}; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190676.4]
  assign notCDom_reduced2AbsSigSum = {reducedVec_orReduceBy2__25,reducedVec_orReduceBy2__24,reducedVec_orReduceBy2__23,reducedVec_orReduceBy2__22,reducedVec_orReduceBy2__21,reducedVec_orReduceBy2__20,reducedVec_orReduceBy2__19,_T_137,_T_132}; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190684.4]
  assign _T_171 = notCDom_reduced2AbsSigSum[1] ? 5'h18 : 5'h19; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190711.4]
  assign _T_172 = notCDom_reduced2AbsSigSum[2] ? 5'h17 : _T_171; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190712.4]
  assign _T_173 = notCDom_reduced2AbsSigSum[3] ? 5'h16 : _T_172; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190713.4]
  assign _T_174 = notCDom_reduced2AbsSigSum[4] ? 5'h15 : _T_173; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190714.4]
  assign _T_175 = notCDom_reduced2AbsSigSum[5] ? 5'h14 : _T_174; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190715.4]
  assign _T_176 = notCDom_reduced2AbsSigSum[6] ? 5'h13 : _T_175; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190716.4]
  assign _T_177 = notCDom_reduced2AbsSigSum[7] ? 5'h12 : _T_176; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190717.4]
  assign _T_178 = notCDom_reduced2AbsSigSum[8] ? 5'h11 : _T_177; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190718.4]
  assign _T_179 = notCDom_reduced2AbsSigSum[9] ? 5'h10 : _T_178; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190719.4]
  assign _T_180 = notCDom_reduced2AbsSigSum[10] ? 5'hf : _T_179; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190720.4]
  assign _T_181 = notCDom_reduced2AbsSigSum[11] ? 5'he : _T_180; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190721.4]
  assign _T_182 = notCDom_reduced2AbsSigSum[12] ? 5'hd : _T_181; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190722.4]
  assign _T_183 = notCDom_reduced2AbsSigSum[13] ? 5'hc : _T_182; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190723.4]
  assign _T_184 = notCDom_reduced2AbsSigSum[14] ? 5'hb : _T_183; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190724.4]
  assign _T_185 = notCDom_reduced2AbsSigSum[15] ? 5'ha : _T_184; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190725.4]
  assign _T_186 = notCDom_reduced2AbsSigSum[16] ? 5'h9 : _T_185; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190726.4]
  assign _T_187 = notCDom_reduced2AbsSigSum[17] ? 5'h8 : _T_186; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190727.4]
  assign _T_188 = notCDom_reduced2AbsSigSum[18] ? 5'h7 : _T_187; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190728.4]
  assign _T_189 = notCDom_reduced2AbsSigSum[19] ? 5'h6 : _T_188; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190729.4]
  assign _T_190 = notCDom_reduced2AbsSigSum[20] ? 5'h5 : _T_189; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190730.4]
  assign _T_191 = notCDom_reduced2AbsSigSum[21] ? 5'h4 : _T_190; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190731.4]
  assign _T_192 = notCDom_reduced2AbsSigSum[22] ? 5'h3 : _T_191; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190732.4]
  assign _T_193 = notCDom_reduced2AbsSigSum[23] ? 5'h2 : _T_192; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190733.4]
  assign _T_194 = notCDom_reduced2AbsSigSum[24] ? 5'h1 : _T_193; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190734.4]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[25] ? 5'h0 : _T_194; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@190735.4]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56:freechips.rocketchip.system.DefaultRV32Config.fir@190736.4]
  assign _T_195 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69:freechips.rocketchip.system.DefaultRV32Config.fir@190737.4]
  assign _GEN_4 = {{3{_T_195[6]}},_T_195}; // @[MulAddRecFN.scala 243:46:freechips.rocketchip.system.DefaultRV32Config.fir@190738.4]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 243:46:freechips.rocketchip.system.DefaultRV32Config.fir@190740.4]
  assign _GEN_5 = {{63'd0}, in_orReduceBy2}; // @[MulAddRecFN.scala 245:27:freechips.rocketchip.system.DefaultRV32Config.fir@190741.4]
  assign _T_198 = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27:freechips.rocketchip.system.DefaultRV32Config.fir@190741.4]
  assign notCDom_mainSig = _T_198[51:23]; // @[MulAddRecFN.scala 245:50:freechips.rocketchip.system.DefaultRV32Config.fir@190742.4]
  assign in_orReduceBy2_1 = notCDom_reduced2AbsSigSum[12:0]; // @[MulAddRecFN.scala 249:39:freechips.rocketchip.system.DefaultRV32Config.fir@190743.4]
  assign reducedVec_orReduceBy2_1_0 = in_orReduceBy2_1[1:0] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190748.4]
  assign reducedVec_orReduceBy2_1_1 = in_orReduceBy2_1[3:2] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190751.4]
  assign reducedVec_orReduceBy2_1_2 = in_orReduceBy2_1[5:4] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190754.4]
  assign reducedVec_orReduceBy2_1_3 = in_orReduceBy2_1[7:6] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190757.4]
  assign reducedVec_orReduceBy2_1_4 = in_orReduceBy2_1[9:8] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190760.4]
  assign reducedVec_orReduceBy2_1_5 = in_orReduceBy2_1[11:10] != 2'h0; // @[primitives.scala 190:54:freechips.rocketchip.system.DefaultRV32Config.fir@190763.4]
  assign reducedVec_orReduceBy2_1_6 = in_orReduceBy2_1[12]; // @[primitives.scala 193:15:freechips.rocketchip.system.DefaultRV32Config.fir@190765.4]
  assign _T_219 = {reducedVec_orReduceBy2_1_6,reducedVec_orReduceBy2_1_5,reducedVec_orReduceBy2_1_4,reducedVec_orReduceBy2_1_3,reducedVec_orReduceBy2_1_2,reducedVec_orReduceBy2_1_1,reducedVec_orReduceBy2_1_0}; // @[primitives.scala 194:20:freechips.rocketchip.system.DefaultRV32Config.fir@190773.4]
  assign in_inv_1 = ~notCDom_normDistReduced2[4:1]; // @[primitives.scala 118:30:freechips.rocketchip.system.DefaultRV32Config.fir@190775.4]
  assign shift_1 = -17'sh10000 >>> in_inv_1; // @[primitives.scala 160:58:freechips.rocketchip.system.DefaultRV32Config.fir@190776.4]
  assign my_lowMask_1_1 = {shift_1[1],shift_1[2],shift_1[3],shift_1[4],shift_1[5],shift_1[6]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190792.4]
  assign _GEN_6 = {{1'd0}, my_lowMask_1_1}; // @[MulAddRecFN.scala 249:78:freechips.rocketchip.system.DefaultRV32Config.fir@190793.4]
  assign _T_236 = _T_219 & _GEN_6; // @[MulAddRecFN.scala 249:78:freechips.rocketchip.system.DefaultRV32Config.fir@190793.4]
  assign notCDom_reduced4SigExtra = _T_236 != 7'h0; // @[MulAddRecFN.scala 251:11:freechips.rocketchip.system.DefaultRV32Config.fir@190794.4]
  assign _T_239 = notCDom_mainSig[2:0] != 3'h0; // @[MulAddRecFN.scala 254:35:freechips.rocketchip.system.DefaultRV32Config.fir@190797.4]
  assign _T_240 = _T_239 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39:freechips.rocketchip.system.DefaultRV32Config.fir@190798.4]
  assign notCDom_sig = {notCDom_mainSig[28:3],_T_240}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190799.4]
  assign notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[MulAddRecFN.scala 257:50:freechips.rocketchip.system.DefaultRV32Config.fir@190801.4]
  assign _T_242 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36:freechips.rocketchip.system.DefaultRV32Config.fir@190802.4]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_242; // @[MulAddRecFN.scala 259:12:freechips.rocketchip.system.DefaultRV32Config.fir@190803.4]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49:freechips.rocketchip.system.DefaultRV32Config.fir@190804.4]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44:freechips.rocketchip.system.DefaultRV32Config.fir@190805.4]
  assign _T_243 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32:freechips.rocketchip.system.DefaultRV32Config.fir@190806.4]
  assign notNaN_addZeros = _T_243 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58:freechips.rocketchip.system.DefaultRV32Config.fir@190807.4]
  assign _T_244 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31:freechips.rocketchip.system.DefaultRV32Config.fir@190808.4]
  assign _T_245 = io_fromPreMul_isSigNaNAny | _T_244; // @[MulAddRecFN.scala 273:35:freechips.rocketchip.system.DefaultRV32Config.fir@190809.4]
  assign _T_246 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32:freechips.rocketchip.system.DefaultRV32Config.fir@190810.4]
  assign _T_247 = _T_245 | _T_246; // @[MulAddRecFN.scala 274:57:freechips.rocketchip.system.DefaultRV32Config.fir@190811.4]
  assign _T_248 = ~io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 276:10:freechips.rocketchip.system.DefaultRV32Config.fir@190812.4]
  assign _T_250 = _T_248 & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36:freechips.rocketchip.system.DefaultRV32Config.fir@190814.4]
  assign _T_251 = _T_250 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61:freechips.rocketchip.system.DefaultRV32Config.fir@190815.4]
  assign _T_252 = _T_251 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35:freechips.rocketchip.system.DefaultRV32Config.fir@190816.4]
  assign _T_255 = ~io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 285:14:freechips.rocketchip.system.DefaultRV32Config.fir@190822.4]
  assign _T_256 = _T_255 & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42:freechips.rocketchip.system.DefaultRV32Config.fir@190823.4]
  assign _T_258 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27:freechips.rocketchip.system.DefaultRV32Config.fir@190826.4]
  assign _T_259 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31:freechips.rocketchip.system.DefaultRV32Config.fir@190827.4]
  assign _T_260 = _T_258 | _T_259; // @[MulAddRecFN.scala 287:54:freechips.rocketchip.system.DefaultRV32Config.fir@190828.4]
  assign _T_261 = ~roundingMode_min; // @[MulAddRecFN.scala 289:29:freechips.rocketchip.system.DefaultRV32Config.fir@190829.4]
  assign _T_262 = notNaN_addZeros & _T_261; // @[MulAddRecFN.scala 289:26:freechips.rocketchip.system.DefaultRV32Config.fir@190830.4]
  assign _T_263 = _T_262 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48:freechips.rocketchip.system.DefaultRV32Config.fir@190831.4]
  assign _T_264 = _T_263 & CDom_sign; // @[MulAddRecFN.scala 290:36:freechips.rocketchip.system.DefaultRV32Config.fir@190832.4]
  assign _T_265 = _T_260 | _T_264; // @[MulAddRecFN.scala 288:43:freechips.rocketchip.system.DefaultRV32Config.fir@190833.4]
  assign _T_266 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26:freechips.rocketchip.system.DefaultRV32Config.fir@190834.4]
  assign _T_267 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37:freechips.rocketchip.system.DefaultRV32Config.fir@190835.4]
  assign _T_268 = _T_266 & _T_267; // @[MulAddRecFN.scala 291:46:freechips.rocketchip.system.DefaultRV32Config.fir@190836.4]
  assign _T_269 = _T_265 | _T_268; // @[MulAddRecFN.scala 290:48:freechips.rocketchip.system.DefaultRV32Config.fir@190837.4]
  assign _T_270 = ~notNaN_isInfOut; // @[MulAddRecFN.scala 293:10:freechips.rocketchip.system.DefaultRV32Config.fir@190838.4]
  assign _T_271 = ~notNaN_addZeros; // @[MulAddRecFN.scala 293:31:freechips.rocketchip.system.DefaultRV32Config.fir@190839.4]
  assign _T_272 = _T_270 & _T_271; // @[MulAddRecFN.scala 293:28:freechips.rocketchip.system.DefaultRV32Config.fir@190840.4]
  assign _T_273 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17:freechips.rocketchip.system.DefaultRV32Config.fir@190841.4]
  assign _T_274 = _T_272 & _T_273; // @[MulAddRecFN.scala 293:49:freechips.rocketchip.system.DefaultRV32Config.fir@190842.4]
  assign io_invalidExc = _T_247 | _T_252; // @[MulAddRecFN.scala 272:19:freechips.rocketchip.system.DefaultRV32Config.fir@190818.4]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21:freechips.rocketchip.system.DefaultRV32Config.fir@190820.4]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21:freechips.rocketchip.system.DefaultRV32Config.fir@190821.4]
  assign io_rawOut_isZero = notNaN_addZeros | _T_256; // @[MulAddRecFN.scala 283:22:freechips.rocketchip.system.DefaultRV32Config.fir@190825.4]
  assign io_rawOut_sign = _T_269 | _T_274; // @[MulAddRecFN.scala 286:20:freechips.rocketchip.system.DefaultRV32Config.fir@190844.4]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20:freechips.rocketchip.system.DefaultRV32Config.fir@190846.4]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19:freechips.rocketchip.system.DefaultRV32Config.fir@190848.4]
endmodule

