`include "include_module.v"
`ifdef __TLB
module TLB( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116715.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116716.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116717.4]
  output        io_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_req_bits_vaddr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_req_bits_passthrough, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_req_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [4:0]  io_req_bits_cmd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_resp_miss, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output [31:0] io_resp_paddr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_resp_pf_ld, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_resp_pf_st, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_resp_ae_ld, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_resp_ae_st, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_resp_ma_ld, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_resp_ma_st, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_resp_cacheable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_sfence_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_sfence_bits_rs1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_sfence_bits_rs2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_sfence_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output        io_ptw_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  output [19:0] io_ptw_req_bits_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_ae, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [53:0] io_ptw_resp_bits_pte_ppn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_pte_d, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_pte_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_pte_g, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_pte_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_pte_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_pte_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_pte_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_pte_v, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_level, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_resp_bits_homogeneous, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_ptbr_mode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_status_debug, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_status_dprv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_status_mxr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_status_sum, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_0_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_pmp_0_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_0_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_0_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_0_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [29:0] io_ptw_pmp_0_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_ptw_pmp_0_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_1_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_pmp_1_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_1_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_1_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_1_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [29:0] io_ptw_pmp_1_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_ptw_pmp_1_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_2_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_pmp_2_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_2_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_2_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_2_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [29:0] io_ptw_pmp_2_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_ptw_pmp_2_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_3_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_pmp_3_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_3_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_3_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_3_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [29:0] io_ptw_pmp_3_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_ptw_pmp_3_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_4_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_pmp_4_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_4_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_4_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_4_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [29:0] io_ptw_pmp_4_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_ptw_pmp_4_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_5_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_pmp_5_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_5_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_5_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_5_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [29:0] io_ptw_pmp_5_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_ptw_pmp_5_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_6_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_pmp_6_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_6_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_6_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_6_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [29:0] io_ptw_pmp_6_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_ptw_pmp_6_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_7_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [1:0]  io_ptw_pmp_7_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_7_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_7_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input         io_ptw_pmp_7_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [29:0] io_ptw_pmp_7_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
  input  [31:0] io_ptw_pmp_7_mask // @[:freechips.rocketchip.system.DefaultRV32Config.fir@116718.4]
);
  wire [19:0] _2_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire [19:0] _2_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire  _2_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
  wire [1:0] pmp_io_prv; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [31:0] pmp_io_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire  pmp_io_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
  wire [19:0] _2_1_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire [19:0] _2_1_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire  _2_1_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
  wire [19:0] _2_2_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire [19:0] _2_2_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire  _2_2_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
  wire [19:0] _2_3_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire [19:0] _2_3_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire  _2_3_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
  wire [19:0] _2_4_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire [19:0] _2_4_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire  _2_4_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
  wire [19:0] _2_5_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire [19:0] _2_5_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire  _2_5_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
  wire [19:0] _2_6_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire [19:0] _2_6_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire  _2_6_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
  wire [19:0] _2_7_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire [19:0] _2_7_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire  _2_7_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
  wire [19:0] _2_8_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire [19:0] _2_8_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire  _2_8_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
  wire [19:0] _2_9_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire [19:0] _2_9_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire  _2_9_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
  wire [19:0] _2_10_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire [19:0] _2_10_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire  _2_10_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
  wire [19:0] _2_11_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire [19:0] _2_11_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire  _2_11_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
  wire [19:0] _2_12_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire [19:0] _2_12_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire  _2_12_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
  wire [19:0] _2_13_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire [19:0] _2_13_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire  _2_13_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
  wire [19:0] _2_14_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire [19:0] _2_14_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire  _2_14_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
  wire [19:0] _2_15_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire [19:0] _2_15_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire  _2_15_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
  wire [19:0] _2_16_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire [19:0] _2_16_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire  _2_16_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
  wire [19:0] _2_17_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire [19:0] _2_17_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire  _2_17_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
  wire [19:0] _2_18_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire [19:0] _2_18_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire  _2_18_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
  wire [19:0] _2_19_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire [19:0] _2_19_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire  _2_19_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
  wire [19:0] _2_20_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire [19:0] _2_20_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire  _2_20_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
  wire [19:0] _2_21_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire [19:0] _2_21_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire  _2_21_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
  wire [19:0] _2_22_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire [19:0] _2_22_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire  _2_22_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
  wire [19:0] _2_23_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire [19:0] _2_23_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire  _2_23_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
  wire [19:0] _2_24_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire [19:0] _2_24_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire  _2_24_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
  wire [19:0] _2_25_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire [19:0] _2_25_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire  _2_25_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
  wire [19:0] _2_26_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire [19:0] _2_26_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire  _2_26_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
  wire [19:0] _2_27_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire [19:0] _2_27_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire  _2_27_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
  wire [19:0] _2_28_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire [19:0] _2_28_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire  _2_28_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
  wire [19:0] _2_29_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire [19:0] _2_29_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire  _2_29_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
  wire [19:0] _2_30_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire [19:0] _2_30_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire  _2_30_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
  wire [19:0] _2_31_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire [19:0] _2_31_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire  _2_31_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
  wire [19:0] _2_32_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire [19:0] _2_32_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire  _2_32_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
  wire [19:0] _2_33_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire [19:0] _2_33_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire  _2_33_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
  wire [19:0] _2_34_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire [19:0] _2_34_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire  _2_34_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
  wire [19:0] _2_35_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire [19:0] _2_35_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire  _2_35_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
  wire [19:0] _2_36_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire [19:0] _2_36_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire  _2_36_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
  wire [19:0] _2_37_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire [19:0] _2_37_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire  _2_37_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
  wire [19:0] _2_38_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire [19:0] _2_38_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  wire  _2_38_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
  reg [19:0] sectored_entries_0_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_0;
  reg [33:0] sectored_entries_0_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_1;
  reg [33:0] sectored_entries_0_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_2;
  reg [33:0] sectored_entries_0_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_3;
  reg [33:0] sectored_entries_0_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_8;
  reg [19:0] sectored_entries_1_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_9;
  reg [33:0] sectored_entries_1_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_10;
  reg [33:0] sectored_entries_1_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_11;
  reg [33:0] sectored_entries_1_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_12;
  reg [33:0] sectored_entries_1_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_13;
  reg  sectored_entries_1_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_14;
  reg  sectored_entries_1_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_15;
  reg  sectored_entries_1_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_16;
  reg  sectored_entries_1_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_17;
  reg [19:0] sectored_entries_2_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_18;
  reg [33:0] sectored_entries_2_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_19;
  reg [33:0] sectored_entries_2_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_20;
  reg [33:0] sectored_entries_2_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_21;
  reg [33:0] sectored_entries_2_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_22;
  reg  sectored_entries_2_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_23;
  reg  sectored_entries_2_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_24;
  reg  sectored_entries_2_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_25;
  reg  sectored_entries_2_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_26;
  reg [19:0] sectored_entries_3_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_27;
  reg [33:0] sectored_entries_3_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_28;
  reg [33:0] sectored_entries_3_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_29;
  reg [33:0] sectored_entries_3_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_30;
  reg [33:0] sectored_entries_3_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_31;
  reg  sectored_entries_3_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_32;
  reg  sectored_entries_3_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_33;
  reg  sectored_entries_3_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_34;
  reg  sectored_entries_3_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_35;
  reg [19:0] sectored_entries_4_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_36;
  reg [33:0] sectored_entries_4_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_37;
  reg [33:0] sectored_entries_4_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_38;
  reg [33:0] sectored_entries_4_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_39;
  reg [33:0] sectored_entries_4_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_40;
  reg  sectored_entries_4_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_41;
  reg  sectored_entries_4_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_42;
  reg  sectored_entries_4_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_43;
  reg  sectored_entries_4_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_44;
  reg [19:0] sectored_entries_5_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_45;
  reg [33:0] sectored_entries_5_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_46;
  reg [33:0] sectored_entries_5_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_47;
  reg [33:0] sectored_entries_5_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_48;
  reg [33:0] sectored_entries_5_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_49;
  reg  sectored_entries_5_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_50;
  reg  sectored_entries_5_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_51;
  reg  sectored_entries_5_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_52;
  reg  sectored_entries_5_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_53;
  reg [19:0] sectored_entries_6_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_54;
  reg [33:0] sectored_entries_6_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_55;
  reg [33:0] sectored_entries_6_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_56;
  reg [33:0] sectored_entries_6_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_57;
  reg [33:0] sectored_entries_6_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_58;
  reg  sectored_entries_6_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_59;
  reg  sectored_entries_6_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_60;
  reg  sectored_entries_6_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_61;
  reg  sectored_entries_6_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_62;
  reg [19:0] sectored_entries_7_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_63;
  reg [33:0] sectored_entries_7_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_64;
  reg [33:0] sectored_entries_7_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_65;
  reg [33:0] sectored_entries_7_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_66;
  reg [33:0] sectored_entries_7_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [63:0] _RAND_67;
  reg  sectored_entries_7_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_68;
  reg  sectored_entries_7_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_69;
  reg  sectored_entries_7_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_70;
  reg  sectored_entries_7_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@116723.4]
  reg [31:0] _RAND_71;
  reg [19:0] superpage_entries_0_tag; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [31:0] _RAND_72;
  reg [33:0] superpage_entries_0_data_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [63:0] _RAND_73;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [31:0] _RAND_74;
  reg [19:0] superpage_entries_1_tag; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [31:0] _RAND_75;
  reg [33:0] superpage_entries_1_data_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [63:0] _RAND_76;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [31:0] _RAND_77;
  reg [19:0] superpage_entries_2_tag; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [31:0] _RAND_78;
  reg [33:0] superpage_entries_2_data_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [63:0] _RAND_79;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [31:0] _RAND_80;
  reg [19:0] superpage_entries_3_tag; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [31:0] _RAND_81;
  reg [33:0] superpage_entries_3_data_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [63:0] _RAND_82;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@116724.4]
  reg [31:0] _RAND_83;
  reg  special_entry_level; // @[TLB.scala 163:56:freechips.rocketchip.system.DefaultRV32Config.fir@116725.4]
  reg [31:0] _RAND_84;
  reg [19:0] special_entry_tag; // @[TLB.scala 163:56:freechips.rocketchip.system.DefaultRV32Config.fir@116725.4]
  reg [31:0] _RAND_85;
  reg [33:0] special_entry_data_0; // @[TLB.scala 163:56:freechips.rocketchip.system.DefaultRV32Config.fir@116725.4]
  reg [63:0] _RAND_86;
  reg  special_entry_valid_0; // @[TLB.scala 163:56:freechips.rocketchip.system.DefaultRV32Config.fir@116725.4]
  reg [31:0] _RAND_87;
  reg [1:0] state; // @[TLB.scala 168:18:freechips.rocketchip.system.DefaultRV32Config.fir@116726.4]
  reg [31:0] _RAND_88;
  reg [19:0] r_refill_tag; // @[TLB.scala 169:25:freechips.rocketchip.system.DefaultRV32Config.fir@116727.4]
  reg [31:0] _RAND_89;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 170:34:freechips.rocketchip.system.DefaultRV32Config.fir@116728.4]
  reg [31:0] _RAND_90;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 171:33:freechips.rocketchip.system.DefaultRV32Config.fir@116729.4]
  reg [31:0] _RAND_91;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 172:32:freechips.rocketchip.system.DefaultRV32Config.fir@116730.4]
  reg [31:0] _RAND_92;
  reg  r_sectored_hit; // @[TLB.scala 173:27:freechips.rocketchip.system.DefaultRV32Config.fir@116731.4]
  reg [31:0] _RAND_93;
  wire  priv_s; // @[TLB.scala 176:20:freechips.rocketchip.system.DefaultRV32Config.fir@116732.4]
  wire  priv_uses_vm; // @[TLB.scala 177:27:freechips.rocketchip.system.DefaultRV32Config.fir@116733.4]
  wire  _T_2; // @[TLB.scala 178:83:freechips.rocketchip.system.DefaultRV32Config.fir@116736.4]
  wire  _T_3; // @[TLB.scala 178:102:freechips.rocketchip.system.DefaultRV32Config.fir@116737.4]
  wire  vm_enabled; // @[TLB.scala 178:99:freechips.rocketchip.system.DefaultRV32Config.fir@116738.4]
  wire [19:0] vpn; // @[TLB.scala 181:30:freechips.rocketchip.system.DefaultRV32Config.fir@116739.4]
  wire [19:0] refill_ppn; // @[TLB.scala 182:44:freechips.rocketchip.system.DefaultRV32Config.fir@116740.4]
  wire  _T_4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@116742.4]
  wire  _T_5; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@116743.4]
  wire  invalidate_refill; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@116744.4]
  wire  _T_21; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@116775.4]
  wire [9:0] _T_24; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@116786.4]
  wire  _T_25; // @[TLB.scala 121:30:freechips.rocketchip.system.DefaultRV32Config.fir@116787.4]
  wire [19:0] _T_27; // @[TLB.scala 122:30:freechips.rocketchip.system.DefaultRV32Config.fir@116789.4]
  wire [19:0] _T_28; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@116790.4]
  wire [9:0] _T_29; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@116791.4]
  wire [19:0] _T_30; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@116792.4]
  wire [19:0] _T_31; // @[TLB.scala 186:123:freechips.rocketchip.system.DefaultRV32Config.fir@116793.4]
  wire [19:0] _T_32; // @[TLB.scala 186:20:freechips.rocketchip.system.DefaultRV32Config.fir@116794.4]
  wire [19:0] mpu_ppn; // @[TLB.scala 185:20:freechips.rocketchip.system.DefaultRV32Config.fir@116795.4]
  wire [11:0] _T_33; // @[TLB.scala 187:52:freechips.rocketchip.system.DefaultRV32Config.fir@116796.4]
  wire [31:0] mpu_physaddr; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@116797.4]
  wire  _T_34; // @[TLB.scala 188:56:freechips.rocketchip.system.DefaultRV32Config.fir@116798.4]
  wire [2:0] _T_36; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@116800.4]
  wire [2:0] mpu_priv; // @[TLB.scala 188:27:freechips.rocketchip.system.DefaultRV32Config.fir@116801.4]
  wire [31:0] _T_37; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116817.4]
  wire [32:0] _T_38; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116818.4]
  wire [32:0] _T_39; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116819.4]
  wire [32:0] _T_40; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116820.4]
  wire  _T_41; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116821.4]
  wire [31:0] _T_42; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116822.4]
  wire [32:0] _T_43; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116823.4]
  wire [32:0] _T_44; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116824.4]
  wire [32:0] _T_45; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116825.4]
  wire  _T_46; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116826.4]
  wire [31:0] _T_47; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116827.4]
  wire [32:0] _T_48; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116828.4]
  wire [32:0] _T_49; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116829.4]
  wire [32:0] _T_50; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116830.4]
  wire  _T_51; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116831.4]
  wire [32:0] _T_53; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116833.4]
  wire [32:0] _T_54; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116834.4]
  wire [32:0] _T_55; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116835.4]
  wire  _T_56; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116836.4]
  wire [31:0] _T_57; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116837.4]
  wire [32:0] _T_58; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116838.4]
  wire [32:0] _T_59; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116839.4]
  wire [32:0] _T_60; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116840.4]
  wire  _T_61; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116841.4]
  wire [31:0] _T_62; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116842.4]
  wire [32:0] _T_63; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116843.4]
  wire [32:0] _T_64; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116844.4]
  wire [32:0] _T_65; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116845.4]
  wire  _T_66; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116846.4]
  wire [31:0] _T_67; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116847.4]
  wire [32:0] _T_68; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116848.4]
  wire [32:0] _T_69; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116849.4]
  wire [32:0] _T_70; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116850.4]
  wire  _T_71; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116851.4]
  wire  _T_73; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116861.4]
  wire  _T_74; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116862.4]
  wire  _T_75; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116863.4]
  wire  _T_76; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116864.4]
  wire  _T_77; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116865.4]
  wire  legal_address; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116866.4]
  wire [32:0] _T_85; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116874.4]
  wire [32:0] _T_86; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116875.4]
  wire  _T_87; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116876.4]
  wire  cacheable; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@116882.4]
  wire [31:0] _T_142; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116934.4]
  wire [32:0] _T_143; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116935.4]
  wire [32:0] _T_144; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116936.4]
  wire [32:0] _T_145; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116937.4]
  wire  _T_146; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116938.4]
  wire [32:0] _T_163; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116955.4]
  wire [32:0] _T_164; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116956.4]
  wire  _T_165; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116957.4]
  wire  _T_172; // @[TLBPermissions.scala 82:66:freechips.rocketchip.system.DefaultRV32Config.fir@116964.4]
  wire  _T_185; // @[TLB.scala 199:39:freechips.rocketchip.system.DefaultRV32Config.fir@116977.4]
  wire  deny_access_to_debug; // @[TLB.scala 199:48:freechips.rocketchip.system.DefaultRV32Config.fir@116983.4]
  wire  _T_197; // @[TLB.scala 200:44:freechips.rocketchip.system.DefaultRV32Config.fir@116990.4]
  wire  _T_198; // @[TLB.scala 200:41:freechips.rocketchip.system.DefaultRV32Config.fir@116991.4]
  wire  prot_r; // @[TLB.scala 200:66:freechips.rocketchip.system.DefaultRV32Config.fir@116992.4]
  wire [32:0] _T_211; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117005.4]
  wire [32:0] _T_212; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117006.4]
  wire  _T_213; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117007.4]
  wire [31:0] _T_214; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@117008.4]
  wire [32:0] _T_215; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@117009.4]
  wire [32:0] _T_216; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117010.4]
  wire [32:0] _T_217; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117011.4]
  wire  _T_218; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117012.4]
  wire  _T_220; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117014.4]
  wire  _T_221; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117015.4]
  wire  _T_231; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@117026.4]
  wire  _T_233; // @[TLB.scala 201:45:freechips.rocketchip.system.DefaultRV32Config.fir@117028.4]
  wire  prot_w; // @[TLB.scala 201:70:freechips.rocketchip.system.DefaultRV32Config.fir@117029.4]
  wire  prot_al; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@117063.4]
  wire [32:0] _T_300; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117100.4]
  wire [32:0] _T_301; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117101.4]
  wire  _T_302; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117102.4]
  wire  _T_313; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117113.4]
  wire  _T_314; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117114.4]
  wire  _T_330; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@117131.4]
  wire  _T_332; // @[TLB.scala 204:40:freechips.rocketchip.system.DefaultRV32Config.fir@117133.4]
  wire  prot_x; // @[TLB.scala 204:65:freechips.rocketchip.system.DefaultRV32Config.fir@117134.4]
  wire [32:0] _T_357; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117159.4]
  wire [32:0] _T_358; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117160.4]
  wire  _T_359; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117161.4]
  wire [32:0] _T_362; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117164.4]
  wire [32:0] _T_363; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117165.4]
  wire  _T_364; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117166.4]
  wire  _T_370; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117172.4]
  wire  _T_371; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117173.4]
  wire  _T_372; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117174.4]
  wire  prot_eff; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@117180.4]
  wire  _T_377; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117181.4]
  wire  _T_378; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117182.4]
  wire  _T_379; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117183.4]
  wire [19:0] _T_380; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117184.4]
  wire [17:0] _T_381; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117185.4]
  wire  _T_382; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117186.4]
  wire  sector_hits_0; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117187.4]
  wire  _T_383; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117188.4]
  wire  _T_384; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117189.4]
  wire  _T_385; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117190.4]
  wire [19:0] _T_386; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117191.4]
  wire [17:0] _T_387; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117192.4]
  wire  _T_388; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117193.4]
  wire  sector_hits_1; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117194.4]
  wire  _T_389; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117195.4]
  wire  _T_390; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117196.4]
  wire  _T_391; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117197.4]
  wire [19:0] _T_392; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117198.4]
  wire [17:0] _T_393; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117199.4]
  wire  _T_394; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117200.4]
  wire  sector_hits_2; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117201.4]
  wire  _T_395; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117202.4]
  wire  _T_396; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117203.4]
  wire  _T_397; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117204.4]
  wire [19:0] _T_398; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117205.4]
  wire [17:0] _T_399; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117206.4]
  wire  _T_400; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117207.4]
  wire  sector_hits_3; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117208.4]
  wire  _T_401; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117209.4]
  wire  _T_402; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117210.4]
  wire  _T_403; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117211.4]
  wire [19:0] _T_404; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117212.4]
  wire [17:0] _T_405; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117213.4]
  wire  _T_406; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117214.4]
  wire  sector_hits_4; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117215.4]
  wire  _T_407; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117216.4]
  wire  _T_408; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117217.4]
  wire  _T_409; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117218.4]
  wire [19:0] _T_410; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117219.4]
  wire [17:0] _T_411; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117220.4]
  wire  _T_412; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117221.4]
  wire  sector_hits_5; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117222.4]
  wire  _T_413; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117223.4]
  wire  _T_414; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117224.4]
  wire  _T_415; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117225.4]
  wire [19:0] _T_416; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117226.4]
  wire [17:0] _T_417; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117227.4]
  wire  _T_418; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117228.4]
  wire  sector_hits_6; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117229.4]
  wire  _T_419; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117230.4]
  wire  _T_420; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117231.4]
  wire  _T_421; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117232.4]
  wire [19:0] _T_422; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117233.4]
  wire [17:0] _T_423; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117234.4]
  wire  _T_424; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117235.4]
  wire  sector_hits_7; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117236.4]
  wire [9:0] _T_427; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117239.4]
  wire [9:0] _T_428; // @[TLB.scala 108:86:freechips.rocketchip.system.DefaultRV32Config.fir@117240.4]
  wire  _T_429; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117241.4]
  wire  superpage_hits_0; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117243.4]
  wire [9:0] _T_435; // @[TLB.scala 108:86:freechips.rocketchip.system.DefaultRV32Config.fir@117247.4]
  wire [9:0] _T_440; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117253.4]
  wire  _T_442; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117255.4]
  wire  superpage_hits_1; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117257.4]
  wire [9:0] _T_453; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117267.4]
  wire  _T_455; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117269.4]
  wire  superpage_hits_2; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117271.4]
  wire [9:0] _T_466; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117281.4]
  wire  _T_468; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117283.4]
  wire  superpage_hits_3; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117285.4]
  wire [1:0] _T_477; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@117293.4]
  wire  _GEN_1; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117297.4]
  wire  _GEN_2; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117297.4]
  wire  _GEN_3; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117297.4]
  wire  _T_481; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117297.4]
  wire  hitsVec_0; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117298.4]
  wire  _GEN_5; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117303.4]
  wire  _GEN_6; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117303.4]
  wire  _GEN_7; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117303.4]
  wire  _T_486; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117303.4]
  wire  hitsVec_1; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117304.4]
  wire  _GEN_9; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117309.4]
  wire  _GEN_10; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117309.4]
  wire  _GEN_11; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117309.4]
  wire  _T_491; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117309.4]
  wire  hitsVec_2; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117310.4]
  wire  _GEN_13; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117315.4]
  wire  _GEN_14; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117315.4]
  wire  _GEN_15; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117315.4]
  wire  _T_496; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117315.4]
  wire  hitsVec_3; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117316.4]
  wire  _GEN_17; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117321.4]
  wire  _GEN_18; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117321.4]
  wire  _GEN_19; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117321.4]
  wire  _T_501; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117321.4]
  wire  hitsVec_4; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117322.4]
  wire  _GEN_21; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117327.4]
  wire  _GEN_22; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117327.4]
  wire  _GEN_23; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117327.4]
  wire  _T_506; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117327.4]
  wire  hitsVec_5; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117328.4]
  wire  _GEN_25; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117333.4]
  wire  _GEN_26; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117333.4]
  wire  _GEN_27; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117333.4]
  wire  _T_511; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117333.4]
  wire  hitsVec_6; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117334.4]
  wire  _GEN_29; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117339.4]
  wire  _GEN_30; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117339.4]
  wire  _GEN_31; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117339.4]
  wire  _T_516; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117339.4]
  wire  hitsVec_7; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117340.4]
  wire  hitsVec_8; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117355.4]
  wire  hitsVec_9; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117370.4]
  wire  hitsVec_10; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117385.4]
  wire  hitsVec_11; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117400.4]
  wire [9:0] _T_575; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117403.4]
  wire  _T_577; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117405.4]
  wire  _T_579; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117407.4]
  wire [9:0] _T_582; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117410.4]
  wire  _T_584; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117412.4]
  wire  _T_585; // @[TLB.scala 108:42:freechips.rocketchip.system.DefaultRV32Config.fir@117413.4]
  wire  _T_586; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117414.4]
  wire  hitsVec_12; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117415.4]
  wire [5:0] _T_591; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117420.4]
  wire [12:0] real_hits; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117427.4]
  wire  _T_598; // @[TLB.scala 211:18:freechips.rocketchip.system.DefaultRV32Config.fir@117428.4]
  wire [13:0] hits; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117429.4]
  wire [33:0] _GEN_33; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117436.4]
  wire [33:0] _GEN_34; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117436.4]
  wire [33:0] _GEN_35; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117436.4]
  wire [33:0] _GEN_37; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117477.4]
  wire [33:0] _GEN_38; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117477.4]
  wire [33:0] _GEN_39; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117477.4]
  wire [33:0] _GEN_41; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117518.4]
  wire [33:0] _GEN_42; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117518.4]
  wire [33:0] _GEN_43; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117518.4]
  wire [33:0] _GEN_45; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117559.4]
  wire [33:0] _GEN_46; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117559.4]
  wire [33:0] _GEN_47; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117559.4]
  wire [33:0] _GEN_49; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117600.4]
  wire [33:0] _GEN_50; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117600.4]
  wire [33:0] _GEN_51; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117600.4]
  wire [33:0] _GEN_53; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117641.4]
  wire [33:0] _GEN_54; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117641.4]
  wire [33:0] _GEN_55; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117641.4]
  wire [33:0] _GEN_57; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117682.4]
  wire [33:0] _GEN_58; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117682.4]
  wire [33:0] _GEN_59; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117682.4]
  wire [33:0] _GEN_61; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117723.4]
  wire [33:0] _GEN_62; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117723.4]
  wire [33:0] _GEN_63; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117723.4]
  wire  _T_758; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@117788.4]
  wire [9:0] _T_761; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117799.4]
  wire [19:0] _T_765; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117803.4]
  wire [9:0] _T_766; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117804.4]
  wire [19:0] _T_767; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117805.4]
  wire  _T_782; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@117835.4]
  wire [9:0] _T_785; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117846.4]
  wire [19:0] _T_789; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117850.4]
  wire [9:0] _T_790; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117851.4]
  wire [19:0] _T_791; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117852.4]
  wire  _T_806; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@117882.4]
  wire [9:0] _T_809; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117893.4]
  wire [19:0] _T_813; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117897.4]
  wire [9:0] _T_814; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117898.4]
  wire [19:0] _T_815; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117899.4]
  wire  _T_830; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@117929.4]
  wire [9:0] _T_833; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117940.4]
  wire [19:0] _T_837; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117944.4]
  wire [9:0] _T_838; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117945.4]
  wire [19:0] _T_839; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117946.4]
  wire [9:0] _T_857; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117987.4]
  wire [19:0] _T_861; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117991.4]
  wire [9:0] _T_862; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117992.4]
  wire [19:0] _T_863; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117993.4]
  wire [19:0] _T_865; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117995.4]
  wire [19:0] _T_866; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117996.4]
  wire [19:0] _T_867; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117997.4]
  wire [19:0] _T_868; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117998.4]
  wire [19:0] _T_869; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117999.4]
  wire [19:0] _T_870; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118000.4]
  wire [19:0] _T_871; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118001.4]
  wire [19:0] _T_872; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118002.4]
  wire [19:0] _T_873; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118003.4]
  wire [19:0] _T_874; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118004.4]
  wire [19:0] _T_875; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118005.4]
  wire [19:0] _T_876; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118006.4]
  wire [19:0] _T_877; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118007.4]
  wire [19:0] _T_878; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118008.4]
  wire [19:0] _T_879; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118009.4]
  wire [19:0] _T_880; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118010.4]
  wire [19:0] _T_881; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118011.4]
  wire [19:0] _T_882; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118012.4]
  wire [19:0] _T_883; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118013.4]
  wire [19:0] _T_884; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118014.4]
  wire [19:0] _T_885; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118015.4]
  wire [19:0] _T_886; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118016.4]
  wire [19:0] _T_887; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118017.4]
  wire [19:0] _T_888; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118018.4]
  wire [19:0] _T_889; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118019.4]
  wire [19:0] _T_890; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118020.4]
  wire [19:0] ppn; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118021.4]
  wire  _T_892; // @[TLB.scala 215:22:freechips.rocketchip.system.DefaultRV32Config.fir@118024.4]
  wire  _T_893; // @[TLB.scala 215:19:freechips.rocketchip.system.DefaultRV32Config.fir@118025.4]
  wire  _T_895; // @[TLB.scala 221:25:freechips.rocketchip.system.DefaultRV32Config.fir@118032.6]
  wire  _T_896; // @[PTW.scala 68:47:freechips.rocketchip.system.DefaultRV32Config.fir@118035.6]
  wire  _T_897; // @[PTW.scala 68:44:freechips.rocketchip.system.DefaultRV32Config.fir@118036.6]
  wire  _T_898; // @[PTW.scala 68:38:freechips.rocketchip.system.DefaultRV32Config.fir@118037.6]
  wire  _T_899; // @[PTW.scala 68:32:freechips.rocketchip.system.DefaultRV32Config.fir@118038.6]
  wire  _T_900; // @[PTW.scala 68:52:freechips.rocketchip.system.DefaultRV32Config.fir@118039.6]
  wire  _T_901; // @[PTW.scala 72:35:freechips.rocketchip.system.DefaultRV32Config.fir@118040.6]
  wire  _T_907; // @[PTW.scala 73:35:freechips.rocketchip.system.DefaultRV32Config.fir@118047.6]
  wire  _T_908; // @[PTW.scala 73:40:freechips.rocketchip.system.DefaultRV32Config.fir@118048.6]
  wire  _T_914; // @[PTW.scala 74:35:freechips.rocketchip.system.DefaultRV32Config.fir@118055.6]
  wire  _T_915; // @[TLB.scala 234:37:freechips.rocketchip.system.DefaultRV32Config.fir@118064.6]
  wire [6:0] _T_923; // @[TLB.scala 136:26:freechips.rocketchip.system.DefaultRV32Config.fir@118076.8]
  wire [33:0] _T_931; // @[TLB.scala 136:26:freechips.rocketchip.system.DefaultRV32Config.fir@118084.8]
  wire  _T_932; // @[TLB.scala 236:40:freechips.rocketchip.system.DefaultRV32Config.fir@118088.8]
  wire  _T_933; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@118090.10]
  wire  _GEN_66; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@118091.10]
  wire  _T_948; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@118111.10]
  wire  _GEN_70; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@118112.10]
  wire  _T_963; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@118132.10]
  wire  _GEN_74; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@118133.10]
  wire  _T_978; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@118153.10]
  wire  _GEN_78; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@118154.10]
  wire [2:0] _T_993; // @[TLB.scala 241:22:freechips.rocketchip.system.DefaultRV32Config.fir@118176.10]
  wire  _T_994; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118177.10]
  wire  _T_995; // @[TLB.scala 243:15:freechips.rocketchip.system.DefaultRV32Config.fir@118179.12]
  wire  _GEN_80; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118180.12]
  wire  _GEN_81; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118180.12]
  wire  _GEN_82; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118180.12]
  wire  _GEN_83; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118180.12]
  wire [1:0] _T_996; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@118188.12]
  wire  _GEN_950; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  wire  _GEN_84; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  wire  _GEN_951; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  wire  _GEN_85; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  wire  _GEN_952; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  wire  _GEN_86; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  wire  _GEN_953; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  wire  _GEN_87; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  wire  _GEN_92; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118178.10]
  wire  _GEN_93; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118178.10]
  wire  _GEN_94; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118178.10]
  wire  _GEN_95; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118178.10]
  wire  _T_1011; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118206.10]
  wire  _GEN_102; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118209.12]
  wire  _GEN_103; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118209.12]
  wire  _GEN_104; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118209.12]
  wire  _GEN_105; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118209.12]
  wire  _GEN_106; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118218.12]
  wire  _GEN_107; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118218.12]
  wire  _GEN_108; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118218.12]
  wire  _GEN_109; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118218.12]
  wire  _GEN_114; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118207.10]
  wire  _GEN_115; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118207.10]
  wire  _GEN_116; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118207.10]
  wire  _GEN_117; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118207.10]
  wire  _T_1028; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118235.10]
  wire  _GEN_124; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118238.12]
  wire  _GEN_125; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118238.12]
  wire  _GEN_126; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118238.12]
  wire  _GEN_127; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118238.12]
  wire  _GEN_128; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118247.12]
  wire  _GEN_129; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118247.12]
  wire  _GEN_130; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118247.12]
  wire  _GEN_131; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118247.12]
  wire  _GEN_136; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118236.10]
  wire  _GEN_137; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118236.10]
  wire  _GEN_138; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118236.10]
  wire  _GEN_139; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118236.10]
  wire  _T_1045; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118264.10]
  wire  _GEN_146; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118267.12]
  wire  _GEN_147; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118267.12]
  wire  _GEN_148; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118267.12]
  wire  _GEN_149; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118267.12]
  wire  _GEN_150; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118276.12]
  wire  _GEN_151; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118276.12]
  wire  _GEN_152; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118276.12]
  wire  _GEN_153; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118276.12]
  wire  _GEN_158; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118265.10]
  wire  _GEN_159; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118265.10]
  wire  _GEN_160; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118265.10]
  wire  _GEN_161; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118265.10]
  wire  _T_1062; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118293.10]
  wire  _GEN_168; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118296.12]
  wire  _GEN_169; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118296.12]
  wire  _GEN_170; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118296.12]
  wire  _GEN_171; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118296.12]
  wire  _GEN_172; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118305.12]
  wire  _GEN_173; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118305.12]
  wire  _GEN_174; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118305.12]
  wire  _GEN_175; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118305.12]
  wire  _GEN_180; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118294.10]
  wire  _GEN_181; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118294.10]
  wire  _GEN_182; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118294.10]
  wire  _GEN_183; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118294.10]
  wire  _T_1079; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118322.10]
  wire  _GEN_190; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118325.12]
  wire  _GEN_191; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118325.12]
  wire  _GEN_192; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118325.12]
  wire  _GEN_193; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118325.12]
  wire  _GEN_194; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118334.12]
  wire  _GEN_195; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118334.12]
  wire  _GEN_196; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118334.12]
  wire  _GEN_197; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118334.12]
  wire  _GEN_202; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118323.10]
  wire  _GEN_203; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118323.10]
  wire  _GEN_204; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118323.10]
  wire  _GEN_205; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118323.10]
  wire  _T_1096; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118351.10]
  wire  _GEN_212; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118354.12]
  wire  _GEN_213; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118354.12]
  wire  _GEN_214; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118354.12]
  wire  _GEN_215; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118354.12]
  wire  _GEN_216; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118363.12]
  wire  _GEN_217; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118363.12]
  wire  _GEN_218; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118363.12]
  wire  _GEN_219; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118363.12]
  wire  _GEN_224; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118352.10]
  wire  _GEN_225; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118352.10]
  wire  _GEN_226; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118352.10]
  wire  _GEN_227; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118352.10]
  wire  _T_1113; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118380.10]
  wire  _GEN_234; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118383.12]
  wire  _GEN_235; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118383.12]
  wire  _GEN_236; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118383.12]
  wire  _GEN_237; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118383.12]
  wire  _GEN_238; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118392.12]
  wire  _GEN_239; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118392.12]
  wire  _GEN_240; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118392.12]
  wire  _GEN_241; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118392.12]
  wire  _GEN_246; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118381.10]
  wire  _GEN_247; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118381.10]
  wire  _GEN_248; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118381.10]
  wire  _GEN_249; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118381.10]
  wire  _GEN_258; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_262; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_266; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_270; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_272; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_273; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_274; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_275; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_282; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_283; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_284; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_285; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_292; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_293; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_294; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_295; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_302; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_303; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_304; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_305; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_312; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_313; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_314; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_315; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_322; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_323; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_324; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_325; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_332; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_333; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_334; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_335; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_342; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_343; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_344; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_345; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  wire  _GEN_354; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_358; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_362; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_366; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_370; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_372; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_373; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_374; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_375; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_382; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_383; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_384; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_385; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_392; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_393; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_394; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_395; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_402; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_403; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_404; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_405; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_412; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_413; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_414; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_415; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_422; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_423; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_424; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_425; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_432; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_433; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_434; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_435; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_442; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_443; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_444; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_445; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  wire  _GEN_454; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_458; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_462; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_466; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_470; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_472; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_473; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_474; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_475; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_482; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_483; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_484; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_485; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_492; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_493; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_494; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_495; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_502; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_503; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_504; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_505; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_512; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_513; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_514; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_515; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_522; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_523; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_524; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_525; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_532; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_533; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_534; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_535; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_542; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_543; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_544; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire  _GEN_545; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  wire [5:0] _T_1575; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119431.4]
  wire [13:0] ptw_ae_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119439.4]
  wire  _T_1583; // @[TLB.scala 253:24:freechips.rocketchip.system.DefaultRV32Config.fir@119440.4]
  wire  _T_1584; // @[TLB.scala 253:32:freechips.rocketchip.system.DefaultRV32Config.fir@119441.4]
  wire [5:0] _T_1589; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119446.4]
  wire [12:0] _T_1596; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119453.4]
  wire [12:0] _T_1597; // @[TLB.scala 253:23:freechips.rocketchip.system.DefaultRV32Config.fir@119454.4]
  wire [12:0] _T_1610; // @[TLB.scala 253:98:freechips.rocketchip.system.DefaultRV32Config.fir@119467.4]
  wire [12:0] _T_1611; // @[TLB.scala 253:89:freechips.rocketchip.system.DefaultRV32Config.fir@119468.4]
  wire [12:0] priv_rw_ok; // @[TLB.scala 253:84:freechips.rocketchip.system.DefaultRV32Config.fir@119469.4]
  wire [5:0] _T_1641; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119500.4]
  wire [12:0] _T_1648; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119507.4]
  wire [5:0] _T_1653; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119512.4]
  wire [12:0] _T_1660; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119519.4]
  wire [12:0] _T_1661; // @[TLB.scala 255:73:freechips.rocketchip.system.DefaultRV32Config.fir@119520.4]
  wire [12:0] _T_1662; // @[TLB.scala 255:68:freechips.rocketchip.system.DefaultRV32Config.fir@119521.4]
  wire [12:0] _T_1663; // @[TLB.scala 255:40:freechips.rocketchip.system.DefaultRV32Config.fir@119522.4]
  wire [13:0] r_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119523.4]
  wire [5:0] _T_1668; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119528.4]
  wire [12:0] _T_1675; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119535.4]
  wire [12:0] _T_1676; // @[TLB.scala 256:40:freechips.rocketchip.system.DefaultRV32Config.fir@119536.4]
  wire [13:0] w_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119537.4]
  wire [1:0] _T_1691; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119553.4]
  wire [5:0] _T_1696; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119558.4]
  wire [13:0] _T_1703; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119565.4]
  wire [13:0] _T_1704; // @[TLB.scala 258:89:freechips.rocketchip.system.DefaultRV32Config.fir@119566.4]
  wire [13:0] pr_array; // @[TLB.scala 258:87:freechips.rocketchip.system.DefaultRV32Config.fir@119567.4]
  wire [1:0] _T_1706; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119569.4]
  wire [5:0] _T_1711; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119574.4]
  wire [13:0] _T_1718; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119581.4]
  wire [13:0] pw_array; // @[TLB.scala 259:87:freechips.rocketchip.system.DefaultRV32Config.fir@119583.4]
  wire [1:0] _T_1736; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119601.4]
  wire [5:0] _T_1741; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119606.4]
  wire [13:0] eff_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119613.4]
  wire [1:0] _T_1749; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119615.4]
  wire [5:0] _T_1754; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119620.4]
  wire [13:0] c_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119627.4]
  wire [1:0] _T_1762; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119629.4]
  wire [5:0] _T_1767; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119634.4]
  wire [13:0] paa_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119641.4]
  wire [5:0] _T_1780; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119648.4]
  wire [13:0] pal_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119655.4]
  wire [13:0] paa_array_if_cached; // @[TLB.scala 265:39:freechips.rocketchip.system.DefaultRV32Config.fir@119657.4]
  wire [13:0] pal_array_if_cached; // @[TLB.scala 266:39:freechips.rocketchip.system.DefaultRV32Config.fir@119659.4]
  wire [3:0] _T_1802; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@119674.4]
  wire [3:0] _T_1804; // @[TLB.scala 269:69:freechips.rocketchip.system.DefaultRV32Config.fir@119676.4]
  wire [31:0] _GEN_982; // @[TLB.scala 269:39:freechips.rocketchip.system.DefaultRV32Config.fir@119677.4]
  wire [31:0] _T_1805; // @[TLB.scala 269:39:freechips.rocketchip.system.DefaultRV32Config.fir@119677.4]
  wire  misaligned; // @[TLB.scala 269:75:freechips.rocketchip.system.DefaultRV32Config.fir@119678.4]
  wire  _T_1806; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119679.4]
  wire  _T_1807; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119680.4]
  wire  cmd_lrsc; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119681.4]
  wire  _T_1809; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119683.4]
  wire  _T_1810; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119684.4]
  wire  _T_1811; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119685.4]
  wire  _T_1812; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119686.4]
  wire  _T_1813; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119687.4]
  wire  _T_1814; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119688.4]
  wire  cmd_amo_logical; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119689.4]
  wire  _T_1816; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119691.4]
  wire  _T_1817; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119692.4]
  wire  _T_1818; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119693.4]
  wire  _T_1819; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119694.4]
  wire  _T_1820; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119695.4]
  wire  _T_1821; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119696.4]
  wire  _T_1822; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119697.4]
  wire  _T_1823; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119698.4]
  wire  cmd_amo_arithmetic; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119699.4]
  wire  _T_1825; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@119701.4]
  wire  _T_1827; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@119703.4]
  wire  _T_1829; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@119705.4]
  wire  _T_1846; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@119722.4]
  wire  cmd_read; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@119723.4]
  wire  _T_1847; // @[Consts.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@119724.4]
  wire  _T_1848; // @[Consts.scala 83:49:freechips.rocketchip.system.DefaultRV32Config.fir@119725.4]
  wire  _T_1849; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@119726.4]
  wire  _T_1851; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@119728.4]
  wire  cmd_write; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@119746.4]
  wire  _T_1869; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119747.4]
  wire  _T_1870; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119748.4]
  wire  _T_1871; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119749.4]
  wire  cmd_write_perms; // @[TLB.scala 285:35:freechips.rocketchip.system.DefaultRV32Config.fir@119750.4]
  wire [13:0] _T_1872; // @[TLB.scala 290:8:freechips.rocketchip.system.DefaultRV32Config.fir@119752.4]
  wire [13:0] _T_1873; // @[TLB.scala 291:19:freechips.rocketchip.system.DefaultRV32Config.fir@119753.4]
  wire [13:0] _T_1874; // @[TLB.scala 291:8:freechips.rocketchip.system.DefaultRV32Config.fir@119754.4]
  wire [13:0] ae_array; // @[TLB.scala 290:37:freechips.rocketchip.system.DefaultRV32Config.fir@119755.4]
  wire [13:0] _T_1875; // @[TLB.scala 292:46:freechips.rocketchip.system.DefaultRV32Config.fir@119756.4]
  wire [13:0] _T_1876; // @[TLB.scala 292:44:freechips.rocketchip.system.DefaultRV32Config.fir@119757.4]
  wire [13:0] ae_ld_array; // @[TLB.scala 292:24:freechips.rocketchip.system.DefaultRV32Config.fir@119758.4]
  wire [13:0] _T_1877; // @[TLB.scala 294:37:freechips.rocketchip.system.DefaultRV32Config.fir@119759.4]
  wire [13:0] _T_1878; // @[TLB.scala 294:35:freechips.rocketchip.system.DefaultRV32Config.fir@119760.4]
  wire [13:0] _T_1879; // @[TLB.scala 294:8:freechips.rocketchip.system.DefaultRV32Config.fir@119761.4]
  wire [13:0] _T_1880; // @[TLB.scala 295:26:freechips.rocketchip.system.DefaultRV32Config.fir@119762.4]
  wire [13:0] _T_1881; // @[TLB.scala 295:8:freechips.rocketchip.system.DefaultRV32Config.fir@119763.4]
  wire [13:0] _T_1882; // @[TLB.scala 294:53:freechips.rocketchip.system.DefaultRV32Config.fir@119764.4]
  wire [13:0] _T_1883; // @[TLB.scala 296:29:freechips.rocketchip.system.DefaultRV32Config.fir@119765.4]
  wire [13:0] _T_1884; // @[TLB.scala 296:8:freechips.rocketchip.system.DefaultRV32Config.fir@119766.4]
  wire [13:0] ae_st_array; // @[TLB.scala 295:53:freechips.rocketchip.system.DefaultRV32Config.fir@119767.4]
  wire  _T_1892; // @[TLB.scala 301:36:freechips.rocketchip.system.DefaultRV32Config.fir@119776.4]
  wire [13:0] _T_1893; // @[TLB.scala 301:49:freechips.rocketchip.system.DefaultRV32Config.fir@119777.4]
  wire [13:0] ma_ld_array; // @[TLB.scala 301:24:freechips.rocketchip.system.DefaultRV32Config.fir@119778.4]
  wire  _T_1894; // @[TLB.scala 302:36:freechips.rocketchip.system.DefaultRV32Config.fir@119779.4]
  wire [13:0] ma_st_array; // @[TLB.scala 302:24:freechips.rocketchip.system.DefaultRV32Config.fir@119781.4]
  wire [13:0] _T_1896; // @[TLB.scala 303:45:freechips.rocketchip.system.DefaultRV32Config.fir@119782.4]
  wire [13:0] _T_1897; // @[TLB.scala 303:35:freechips.rocketchip.system.DefaultRV32Config.fir@119783.4]
  wire [13:0] pf_ld_array; // @[TLB.scala 303:24:freechips.rocketchip.system.DefaultRV32Config.fir@119784.4]
  wire [13:0] _T_1898; // @[TLB.scala 304:52:freechips.rocketchip.system.DefaultRV32Config.fir@119785.4]
  wire [13:0] _T_1899; // @[TLB.scala 304:42:freechips.rocketchip.system.DefaultRV32Config.fir@119786.4]
  wire [13:0] pf_st_array; // @[TLB.scala 304:24:freechips.rocketchip.system.DefaultRV32Config.fir@119787.4]
  wire  tlb_hit; // @[TLB.scala 307:27:freechips.rocketchip.system.DefaultRV32Config.fir@119790.4]
  wire  _T_1903; // @[TLB.scala 308:43:freechips.rocketchip.system.DefaultRV32Config.fir@119793.4]
  wire  tlb_miss; // @[TLB.scala 308:40:freechips.rocketchip.system.DefaultRV32Config.fir@119794.4]
  reg [6:0] _T_1904; // @[Replacement.scala 41:30:freechips.rocketchip.system.DefaultRV32Config.fir@119795.4]
  reg [31:0] _RAND_94;
  reg [2:0] _T_1905; // @[Replacement.scala 41:30:freechips.rocketchip.system.DefaultRV32Config.fir@119796.4]
  reg [31:0] _RAND_95;
  wire  _T_1906; // @[TLB.scala 312:22:freechips.rocketchip.system.DefaultRV32Config.fir@119797.4]
  wire  _T_1907; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119799.6]
  wire  _T_1908; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119800.6]
  wire  _T_1909; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119801.6]
  wire  _T_1910; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119802.6]
  wire  _T_1911; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119803.6]
  wire  _T_1912; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119804.6]
  wire  _T_1913; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119805.6]
  wire [7:0] _T_1920; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119813.8]
  wire [3:0] _T_1921; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@119814.8]
  wire [3:0] _T_1922; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@119815.8]
  wire  _T_1923; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@119816.8]
  wire [3:0] _T_1924; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@119817.8]
  wire [1:0] _T_1925; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@119818.8]
  wire [1:0] _T_1926; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@119819.8]
  wire  _T_1927; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@119820.8]
  wire [1:0] _T_1928; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@119821.8]
  wire  _T_1929; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@119822.8]
  wire [2:0] _T_1931; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119824.8]
  wire [7:0] _T_1932; // @[Replacement.scala 46:28:freechips.rocketchip.system.DefaultRV32Config.fir@119825.8]
  wire  _T_1933; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119826.8]
  wire  _T_1934; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119827.8]
  wire [7:0] _T_1936; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119829.8]
  wire [7:0] _T_1937; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119830.8]
  wire [7:0] _T_1938; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119831.8]
  wire [7:0] _T_1939; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119832.8]
  wire [7:0] _T_1940; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119833.8]
  wire [1:0] _T_1941; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119834.8]
  wire  _T_1942; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119835.8]
  wire  _T_1943; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119836.8]
  wire [3:0] _T_1944; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119837.8]
  wire [7:0] _GEN_983; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119838.8]
  wire [7:0] _T_1945; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119838.8]
  wire [7:0] _T_1946; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119839.8]
  wire [7:0] _T_1947; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119840.8]
  wire [7:0] _T_1948; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119841.8]
  wire [7:0] _T_1949; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119842.8]
  wire [2:0] _T_1950; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119843.8]
  wire  _T_1951; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119844.8]
  wire  _T_1952; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119845.8]
  wire [7:0] _T_1953; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119846.8]
  wire [7:0] _T_1954; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119847.8]
  wire [7:0] _T_1955; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119848.8]
  wire [7:0] _T_1956; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119849.8]
  wire [7:0] _T_1957; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119850.8]
  wire [7:0] _T_1958; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119851.8]
  wire [6:0] _T_1960; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@119853.8]
  wire  _T_1961; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119856.6]
  wire  _T_1962; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119857.6]
  wire  _T_1963; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119858.6]
  wire [3:0] _T_1966; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119862.8]
  wire [1:0] _T_1967; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@119863.8]
  wire [1:0] _T_1968; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@119864.8]
  wire  _T_1969; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@119865.8]
  wire [1:0] _T_1970; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@119866.8]
  wire  _T_1971; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@119867.8]
  wire [1:0] _T_1972; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119868.8]
  wire [3:0] _T_1973; // @[Replacement.scala 46:28:freechips.rocketchip.system.DefaultRV32Config.fir@119869.8]
  wire  _T_1974; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119870.8]
  wire  _T_1975; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119871.8]
  wire [3:0] _T_1977; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119873.8]
  wire [3:0] _T_1978; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119874.8]
  wire [3:0] _T_1979; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119875.8]
  wire [3:0] _T_1980; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119876.8]
  wire [3:0] _T_1981; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119877.8]
  wire [1:0] _T_1982; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119878.8]
  wire  _T_1983; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119879.8]
  wire  _T_1984; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119880.8]
  wire [3:0] _T_1985; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119881.8]
  wire [3:0] _T_1986; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119882.8]
  wire [3:0] _T_1987; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119883.8]
  wire [3:0] _T_1988; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119884.8]
  wire [3:0] _T_1989; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119885.8]
  wire [3:0] _T_1990; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119886.8]
  wire [2:0] _T_1992; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@119888.8]
  wire [5:0] _T_1993; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119892.4]
  wire [2:0] _T_1994; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119893.4]
  wire  _T_1995; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119894.4]
  wire [1:0] _T_1997; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119896.4]
  wire  _T_1998; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119897.4]
  wire  _T_2000; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119899.4]
  wire  _T_2002; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119901.4]
  wire  _T_2004; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119903.4]
  wire  _T_2006; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119905.4]
  wire  _T_2008; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119907.4]
  wire  _T_2009; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119908.4]
  wire [2:0] _T_2010; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119909.4]
  wire  _T_2011; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119910.4]
  wire [1:0] _T_2013; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119912.4]
  wire  _T_2014; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119913.4]
  wire  _T_2016; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119915.4]
  wire  _T_2018; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119917.4]
  wire  _T_2020; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119919.4]
  wire  _T_2022; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119921.4]
  wire  _T_2024; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119923.4]
  wire  _T_2025; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119924.4]
  wire  _T_2026; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119925.4]
  wire  _T_2027; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@119926.4]
  wire  _T_2028; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119927.4]
  wire  _T_2029; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119928.4]
  wire [6:0] _T_2030; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119929.4]
  wire [2:0] _T_2031; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119930.4]
  wire  _T_2032; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119931.4]
  wire [1:0] _T_2034; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119933.4]
  wire  _T_2035; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119934.4]
  wire  _T_2037; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119936.4]
  wire  _T_2039; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119938.4]
  wire  _T_2041; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119940.4]
  wire  _T_2043; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119942.4]
  wire  _T_2045; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119944.4]
  wire  _T_2046; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119945.4]
  wire [3:0] _T_2047; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119946.4]
  wire [1:0] _T_2048; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119947.4]
  wire  _T_2049; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119948.4]
  wire  _T_2051; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119950.4]
  wire  _T_2053; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119952.4]
  wire  _T_2055; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119954.4]
  wire [1:0] _T_2057; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119956.4]
  wire  _T_2058; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119957.4]
  wire  _T_2060; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119959.4]
  wire  _T_2062; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119961.4]
  wire  _T_2064; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119963.4]
  wire  _T_2066; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119965.4]
  wire  _T_2067; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@119966.4]
  wire  _T_2068; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119967.4]
  wire  _T_2069; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119968.4]
  wire  _T_2070; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119969.4]
  wire  _T_2071; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@119970.4]
  wire  _T_2072; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119971.4]
  wire  _T_2073; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119972.4]
  wire  _T_2075; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@119974.4]
  wire  _T_2076; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119975.4]
  wire  multipleHits; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119976.4]
  wire [13:0] _T_2079; // @[TLB.scala 325:57:freechips.rocketchip.system.DefaultRV32Config.fir@119980.4]
  wire [13:0] _T_2083; // @[TLB.scala 326:64:freechips.rocketchip.system.DefaultRV32Config.fir@119985.4]
  wire [13:0] _T_2089; // @[TLB.scala 328:33:freechips.rocketchip.system.DefaultRV32Config.fir@119993.4]
  wire [13:0] _T_2091; // @[TLB.scala 329:33:freechips.rocketchip.system.DefaultRV32Config.fir@119996.4]
  wire [13:0] _T_2096; // @[TLB.scala 331:33:freechips.rocketchip.system.DefaultRV32Config.fir@120003.4]
  wire [13:0] _T_2098; // @[TLB.scala 332:33:freechips.rocketchip.system.DefaultRV32Config.fir@120006.4]
  wire [13:0] _T_2100; // @[TLB.scala 334:33:freechips.rocketchip.system.DefaultRV32Config.fir@120010.4]
  wire  _T_2107; // @[TLB.scala 337:29:freechips.rocketchip.system.DefaultRV32Config.fir@120020.4]
  wire  _T_2113; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@120031.4]
  wire  _T_2114; // @[TLB.scala 346:25:freechips.rocketchip.system.DefaultRV32Config.fir@120032.4]
  wire [2:0] _GEN_985; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120040.6]
  wire [3:0] _T_2119; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120040.6]
  wire  _T_2120; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120041.6]
  wire [1:0] _T_2122; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120043.6]
  wire [3:0] _T_2126; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120047.6]
  wire  _T_2127; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120048.6]
  wire [2:0] _T_2129; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120050.6]
  wire [1:0] _T_2130; // @[Replacement.scala 63:8:freechips.rocketchip.system.DefaultRV32Config.fir@120051.6]
  wire [3:0] _T_2133; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120054.6]
  wire  _T_2134; // @[TLB.scala 394:16:freechips.rocketchip.system.DefaultRV32Config.fir@120055.6]
  wire [3:0] _T_2135; // @[TLB.scala 394:43:freechips.rocketchip.system.DefaultRV32Config.fir@120056.6]
  wire  _T_2136; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120057.6]
  wire  _T_2137; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120058.6]
  wire  _T_2138; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120059.6]
  wire [6:0] _GEN_986; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120070.6]
  wire [7:0] _T_2148; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120070.6]
  wire  _T_2149; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120071.6]
  wire [1:0] _T_2151; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120073.6]
  wire [7:0] _T_2155; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120077.6]
  wire  _T_2156; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120078.6]
  wire [2:0] _T_2158; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120080.6]
  wire [7:0] _T_2162; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120084.6]
  wire  _T_2163; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120085.6]
  wire [3:0] _T_2165; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120087.6]
  wire [2:0] _T_2166; // @[Replacement.scala 63:8:freechips.rocketchip.system.DefaultRV32Config.fir@120088.6]
  wire [7:0] _T_2197; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120119.6]
  wire  _T_2198; // @[TLB.scala 394:16:freechips.rocketchip.system.DefaultRV32Config.fir@120120.6]
  wire [7:0] _T_2199; // @[TLB.scala 394:43:freechips.rocketchip.system.DefaultRV32Config.fir@120121.6]
  wire  _T_2200; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120122.6]
  wire  _T_2201; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120123.6]
  wire  _T_2202; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120124.6]
  wire  _T_2203; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120125.6]
  wire  _T_2204; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120126.6]
  wire  _T_2205; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120127.6]
  wire  _T_2206; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120128.6]
  wire  _T_2243; // @[TLB.scala 360:17:freechips.rocketchip.system.DefaultRV32Config.fir@120180.4]
  wire  _T_2244; // @[TLB.scala 360:28:freechips.rocketchip.system.DefaultRV32Config.fir@120181.4]
  wire  _T_2245; // @[TLB.scala 368:14:freechips.rocketchip.system.DefaultRV32Config.fir@120189.6]
  wire [19:0] _T_2246; // @[TLB.scala 368:58:freechips.rocketchip.system.DefaultRV32Config.fir@120190.6]
  wire  _T_2247; // @[TLB.scala 368:72:freechips.rocketchip.system.DefaultRV32Config.fir@120191.6]
  wire  _T_2248; // @[TLB.scala 368:34:freechips.rocketchip.system.DefaultRV32Config.fir@120192.6]
  wire  _T_2250; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@120194.6]
  wire  _T_2251; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@120195.6]
  wire [9:0] _T_2257; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@120209.8]
  wire  _T_2258; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@120210.8]
  wire  _T_2261; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120217.10]
  wire  _T_2273; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120241.10]
  wire  _T_2278; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120252.10]
  wire  _T_2290; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120276.10]
  wire  _T_2295; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120287.10]
  wire  _T_2307; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120311.10]
  wire  _T_2312; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120322.10]
  wire  _T_2324; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120346.10]
  wire  _T_2395; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120508.10]
  wire  _GEN_648; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120509.10]
  wire  _T_2396; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120512.10]
  wire  _GEN_649; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120513.10]
  wire  _T_2397; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120516.10]
  wire  _GEN_650; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120517.10]
  wire  _T_2398; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120520.10]
  wire  _GEN_651; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120521.10]
  wire  _GEN_652; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120367.8]
  wire  _GEN_653; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120367.8]
  wire  _GEN_654; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120367.8]
  wire  _GEN_655; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120367.8]
  wire [9:0] _T_2404; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@120540.8]
  wire  _T_2405; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@120541.8]
  wire  _T_2408; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120548.10]
  wire  _T_2420; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120572.10]
  wire  _T_2425; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120583.10]
  wire  _T_2437; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120607.10]
  wire  _T_2442; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120618.10]
  wire  _T_2454; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120642.10]
  wire  _T_2459; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120653.10]
  wire  _T_2471; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120677.10]
  wire  _T_2542; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120839.10]
  wire  _GEN_676; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120840.10]
  wire  _T_2543; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120843.10]
  wire  _GEN_677; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120844.10]
  wire  _T_2544; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120847.10]
  wire  _GEN_678; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120848.10]
  wire  _T_2545; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120851.10]
  wire  _GEN_679; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120852.10]
  wire  _GEN_680; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120698.8]
  wire  _GEN_681; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120698.8]
  wire  _GEN_682; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120698.8]
  wire  _GEN_683; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120698.8]
  wire [9:0] _T_2551; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@120871.8]
  wire  _T_2552; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@120872.8]
  wire  _T_2555; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120879.10]
  wire  _T_2567; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120903.10]
  wire  _T_2572; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120914.10]
  wire  _T_2584; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120938.10]
  wire  _T_2589; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120949.10]
  wire  _T_2601; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120973.10]
  wire  _T_2606; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120984.10]
  wire  _T_2618; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121008.10]
  wire  _T_2689; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121170.10]
  wire  _GEN_704; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121171.10]
  wire  _T_2690; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121174.10]
  wire  _GEN_705; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121175.10]
  wire  _T_2691; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121178.10]
  wire  _GEN_706; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121179.10]
  wire  _T_2692; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121182.10]
  wire  _GEN_707; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121183.10]
  wire  _GEN_708; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121029.8]
  wire  _GEN_709; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121029.8]
  wire  _GEN_710; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121029.8]
  wire  _GEN_711; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121029.8]
  wire [9:0] _T_2698; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@121202.8]
  wire  _T_2699; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@121203.8]
  wire  _T_2702; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121210.10]
  wire  _T_2714; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121234.10]
  wire  _T_2719; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121245.10]
  wire  _T_2731; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121269.10]
  wire  _T_2736; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121280.10]
  wire  _T_2748; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121304.10]
  wire  _T_2753; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121315.10]
  wire  _T_2765; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121339.10]
  wire  _T_2836; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121501.10]
  wire  _GEN_732; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121502.10]
  wire  _T_2837; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121505.10]
  wire  _GEN_733; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121506.10]
  wire  _T_2838; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121509.10]
  wire  _GEN_734; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121510.10]
  wire  _T_2839; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121513.10]
  wire  _GEN_735; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121514.10]
  wire  _GEN_736; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121360.8]
  wire  _GEN_737; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121360.8]
  wire  _GEN_738; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121360.8]
  wire  _GEN_739; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121360.8]
  wire [9:0] _T_2845; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@121533.8]
  wire  _T_2846; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@121534.8]
  wire  _T_2849; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121541.10]
  wire  _T_2861; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121565.10]
  wire  _T_2866; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121576.10]
  wire  _T_2878; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121600.10]
  wire  _T_2883; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121611.10]
  wire  _T_2895; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121635.10]
  wire  _T_2900; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121646.10]
  wire  _T_2912; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121670.10]
  wire  _T_2983; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121832.10]
  wire  _GEN_760; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121833.10]
  wire  _T_2984; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121836.10]
  wire  _GEN_761; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121837.10]
  wire  _T_2985; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121840.10]
  wire  _GEN_762; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121841.10]
  wire  _T_2986; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121844.10]
  wire  _GEN_763; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121845.10]
  wire  _GEN_764; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121691.8]
  wire  _GEN_765; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121691.8]
  wire  _GEN_766; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121691.8]
  wire  _GEN_767; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121691.8]
  wire [9:0] _T_2992; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@121864.8]
  wire  _T_2993; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@121865.8]
  wire  _T_2996; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121872.10]
  wire  _T_3008; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121896.10]
  wire  _T_3013; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121907.10]
  wire  _T_3025; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121931.10]
  wire  _T_3030; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121942.10]
  wire  _T_3042; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121966.10]
  wire  _T_3047; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121977.10]
  wire  _T_3059; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122001.10]
  wire  _T_3130; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122163.10]
  wire  _GEN_788; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122164.10]
  wire  _T_3131; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122167.10]
  wire  _GEN_789; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122168.10]
  wire  _T_3132; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122171.10]
  wire  _GEN_790; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122172.10]
  wire  _T_3133; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122175.10]
  wire  _GEN_791; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122176.10]
  wire  _GEN_792; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122022.8]
  wire  _GEN_793; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122022.8]
  wire  _GEN_794; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122022.8]
  wire  _GEN_795; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122022.8]
  wire [9:0] _T_3139; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@122195.8]
  wire  _T_3140; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@122196.8]
  wire  _T_3143; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122203.10]
  wire  _T_3155; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122227.10]
  wire  _T_3160; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122238.10]
  wire  _T_3172; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122262.10]
  wire  _T_3177; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122273.10]
  wire  _T_3189; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122297.10]
  wire  _T_3194; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122308.10]
  wire  _T_3206; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122332.10]
  wire  _T_3277; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122494.10]
  wire  _GEN_816; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122495.10]
  wire  _T_3278; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122498.10]
  wire  _GEN_817; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122499.10]
  wire  _T_3279; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122502.10]
  wire  _GEN_818; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122503.10]
  wire  _T_3280; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122506.10]
  wire  _GEN_819; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122507.10]
  wire  _GEN_820; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122353.8]
  wire  _GEN_821; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122353.8]
  wire  _GEN_822; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122353.8]
  wire  _GEN_823; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122353.8]
  wire [9:0] _T_3286; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@122526.8]
  wire  _T_3287; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@122527.8]
  wire  _T_3290; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122534.10]
  wire  _T_3302; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122558.10]
  wire  _T_3307; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122569.10]
  wire  _T_3319; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122593.10]
  wire  _T_3324; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122604.10]
  wire  _T_3336; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122628.10]
  wire  _T_3341; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122639.10]
  wire  _T_3353; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122663.10]
  wire  _T_3424; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122825.10]
  wire  _GEN_844; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122826.10]
  wire  _T_3425; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122829.10]
  wire  _GEN_845; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122830.10]
  wire  _T_3426; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122833.10]
  wire  _GEN_846; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122834.10]
  wire  _T_3427; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122837.10]
  wire  _GEN_847; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122838.10]
  wire  _GEN_848; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122684.8]
  wire  _GEN_849; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122684.8]
  wire  _GEN_850; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122684.8]
  wire  _GEN_851; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122684.8]
  wire  _T_3459; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122904.10]
  wire  _GEN_857; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122905.10]
  wire  _GEN_858; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122868.8]
  wire  _T_3491; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122968.10]
  wire  _GEN_861; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122969.10]
  wire  _GEN_862; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122932.8]
  wire  _T_3523; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@123032.10]
  wire  _GEN_865; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@123033.10]
  wire  _GEN_866; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122996.8]
  wire  _T_3555; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@123096.10]
  wire  _GEN_869; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@123097.10]
  wire  _GEN_870; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@123060.8]
  wire  _T_3587; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@123160.10]
  wire  _GEN_873; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@123161.10]
  wire  _GEN_874; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@123124.8]
  wire  _T_3589; // @[TLB.scala 375:24:freechips.rocketchip.system.DefaultRV32Config.fir@123170.4]
  _2_1 _2 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@116781.4]
    .io_x_ppn(_2_io_x_ppn),
    .io_x_u(_2_io_x_u),
    .io_x_ae(_2_io_x_ae),
    .io_x_sw(_2_io_x_sw),
    .io_x_sx(_2_io_x_sx),
    .io_x_sr(_2_io_x_sr),
    .io_x_pw(_2_io_x_pw),
    .io_x_px(_2_io_x_px),
    .io_x_pr(_2_io_x_pr),
    .io_x_pal(_2_io_x_pal),
    .io_x_paa(_2_io_x_paa),
    .io_x_eff(_2_io_x_eff),
    .io_x_c(_2_io_x_c),
    .io_y_ppn(_2_io_y_ppn),
    .io_y_u(_2_io_y_u),
    .io_y_ae(_2_io_y_ae),
    .io_y_sw(_2_io_y_sw),
    .io_y_sx(_2_io_y_sx),
    .io_y_sr(_2_io_y_sr),
    .io_y_pw(_2_io_y_pw),
    .io_y_px(_2_io_y_px),
    .io_y_pr(_2_io_y_pr),
    .io_y_pal(_2_io_y_pal),
    .io_y_paa(_2_io_y_paa),
    .io_y_eff(_2_io_y_eff),
    .io_y_c(_2_io_y_c)
  );
  PMPChecker pmp ( // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@116802.4]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x)
  );
  _2_1 _2_1 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117467.4]
    .io_x_ppn(_2_1_io_x_ppn),
    .io_x_u(_2_1_io_x_u),
    .io_x_ae(_2_1_io_x_ae),
    .io_x_sw(_2_1_io_x_sw),
    .io_x_sx(_2_1_io_x_sx),
    .io_x_sr(_2_1_io_x_sr),
    .io_x_pw(_2_1_io_x_pw),
    .io_x_px(_2_1_io_x_px),
    .io_x_pr(_2_1_io_x_pr),
    .io_x_pal(_2_1_io_x_pal),
    .io_x_paa(_2_1_io_x_paa),
    .io_x_eff(_2_1_io_x_eff),
    .io_x_c(_2_1_io_x_c),
    .io_y_ppn(_2_1_io_y_ppn),
    .io_y_u(_2_1_io_y_u),
    .io_y_ae(_2_1_io_y_ae),
    .io_y_sw(_2_1_io_y_sw),
    .io_y_sx(_2_1_io_y_sx),
    .io_y_sr(_2_1_io_y_sr),
    .io_y_pw(_2_1_io_y_pw),
    .io_y_px(_2_1_io_y_px),
    .io_y_pr(_2_1_io_y_pr),
    .io_y_pal(_2_1_io_y_pal),
    .io_y_paa(_2_1_io_y_paa),
    .io_y_eff(_2_1_io_y_eff),
    .io_y_c(_2_1_io_y_c)
  );
  _2_1 _2_2 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117508.4]
    .io_x_ppn(_2_2_io_x_ppn),
    .io_x_u(_2_2_io_x_u),
    .io_x_ae(_2_2_io_x_ae),
    .io_x_sw(_2_2_io_x_sw),
    .io_x_sx(_2_2_io_x_sx),
    .io_x_sr(_2_2_io_x_sr),
    .io_x_pw(_2_2_io_x_pw),
    .io_x_px(_2_2_io_x_px),
    .io_x_pr(_2_2_io_x_pr),
    .io_x_pal(_2_2_io_x_pal),
    .io_x_paa(_2_2_io_x_paa),
    .io_x_eff(_2_2_io_x_eff),
    .io_x_c(_2_2_io_x_c),
    .io_y_ppn(_2_2_io_y_ppn),
    .io_y_u(_2_2_io_y_u),
    .io_y_ae(_2_2_io_y_ae),
    .io_y_sw(_2_2_io_y_sw),
    .io_y_sx(_2_2_io_y_sx),
    .io_y_sr(_2_2_io_y_sr),
    .io_y_pw(_2_2_io_y_pw),
    .io_y_px(_2_2_io_y_px),
    .io_y_pr(_2_2_io_y_pr),
    .io_y_pal(_2_2_io_y_pal),
    .io_y_paa(_2_2_io_y_paa),
    .io_y_eff(_2_2_io_y_eff),
    .io_y_c(_2_2_io_y_c)
  );
  _2_1 _2_3 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117549.4]
    .io_x_ppn(_2_3_io_x_ppn),
    .io_x_u(_2_3_io_x_u),
    .io_x_ae(_2_3_io_x_ae),
    .io_x_sw(_2_3_io_x_sw),
    .io_x_sx(_2_3_io_x_sx),
    .io_x_sr(_2_3_io_x_sr),
    .io_x_pw(_2_3_io_x_pw),
    .io_x_px(_2_3_io_x_px),
    .io_x_pr(_2_3_io_x_pr),
    .io_x_pal(_2_3_io_x_pal),
    .io_x_paa(_2_3_io_x_paa),
    .io_x_eff(_2_3_io_x_eff),
    .io_x_c(_2_3_io_x_c),
    .io_y_ppn(_2_3_io_y_ppn),
    .io_y_u(_2_3_io_y_u),
    .io_y_ae(_2_3_io_y_ae),
    .io_y_sw(_2_3_io_y_sw),
    .io_y_sx(_2_3_io_y_sx),
    .io_y_sr(_2_3_io_y_sr),
    .io_y_pw(_2_3_io_y_pw),
    .io_y_px(_2_3_io_y_px),
    .io_y_pr(_2_3_io_y_pr),
    .io_y_pal(_2_3_io_y_pal),
    .io_y_paa(_2_3_io_y_paa),
    .io_y_eff(_2_3_io_y_eff),
    .io_y_c(_2_3_io_y_c)
  );
  _2_1 _2_4 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117590.4]
    .io_x_ppn(_2_4_io_x_ppn),
    .io_x_u(_2_4_io_x_u),
    .io_x_ae(_2_4_io_x_ae),
    .io_x_sw(_2_4_io_x_sw),
    .io_x_sx(_2_4_io_x_sx),
    .io_x_sr(_2_4_io_x_sr),
    .io_x_pw(_2_4_io_x_pw),
    .io_x_px(_2_4_io_x_px),
    .io_x_pr(_2_4_io_x_pr),
    .io_x_pal(_2_4_io_x_pal),
    .io_x_paa(_2_4_io_x_paa),
    .io_x_eff(_2_4_io_x_eff),
    .io_x_c(_2_4_io_x_c),
    .io_y_ppn(_2_4_io_y_ppn),
    .io_y_u(_2_4_io_y_u),
    .io_y_ae(_2_4_io_y_ae),
    .io_y_sw(_2_4_io_y_sw),
    .io_y_sx(_2_4_io_y_sx),
    .io_y_sr(_2_4_io_y_sr),
    .io_y_pw(_2_4_io_y_pw),
    .io_y_px(_2_4_io_y_px),
    .io_y_pr(_2_4_io_y_pr),
    .io_y_pal(_2_4_io_y_pal),
    .io_y_paa(_2_4_io_y_paa),
    .io_y_eff(_2_4_io_y_eff),
    .io_y_c(_2_4_io_y_c)
  );
  _2_1 _2_5 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117631.4]
    .io_x_ppn(_2_5_io_x_ppn),
    .io_x_u(_2_5_io_x_u),
    .io_x_ae(_2_5_io_x_ae),
    .io_x_sw(_2_5_io_x_sw),
    .io_x_sx(_2_5_io_x_sx),
    .io_x_sr(_2_5_io_x_sr),
    .io_x_pw(_2_5_io_x_pw),
    .io_x_px(_2_5_io_x_px),
    .io_x_pr(_2_5_io_x_pr),
    .io_x_pal(_2_5_io_x_pal),
    .io_x_paa(_2_5_io_x_paa),
    .io_x_eff(_2_5_io_x_eff),
    .io_x_c(_2_5_io_x_c),
    .io_y_ppn(_2_5_io_y_ppn),
    .io_y_u(_2_5_io_y_u),
    .io_y_ae(_2_5_io_y_ae),
    .io_y_sw(_2_5_io_y_sw),
    .io_y_sx(_2_5_io_y_sx),
    .io_y_sr(_2_5_io_y_sr),
    .io_y_pw(_2_5_io_y_pw),
    .io_y_px(_2_5_io_y_px),
    .io_y_pr(_2_5_io_y_pr),
    .io_y_pal(_2_5_io_y_pal),
    .io_y_paa(_2_5_io_y_paa),
    .io_y_eff(_2_5_io_y_eff),
    .io_y_c(_2_5_io_y_c)
  );
  _2_1 _2_6 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117672.4]
    .io_x_ppn(_2_6_io_x_ppn),
    .io_x_u(_2_6_io_x_u),
    .io_x_ae(_2_6_io_x_ae),
    .io_x_sw(_2_6_io_x_sw),
    .io_x_sx(_2_6_io_x_sx),
    .io_x_sr(_2_6_io_x_sr),
    .io_x_pw(_2_6_io_x_pw),
    .io_x_px(_2_6_io_x_px),
    .io_x_pr(_2_6_io_x_pr),
    .io_x_pal(_2_6_io_x_pal),
    .io_x_paa(_2_6_io_x_paa),
    .io_x_eff(_2_6_io_x_eff),
    .io_x_c(_2_6_io_x_c),
    .io_y_ppn(_2_6_io_y_ppn),
    .io_y_u(_2_6_io_y_u),
    .io_y_ae(_2_6_io_y_ae),
    .io_y_sw(_2_6_io_y_sw),
    .io_y_sx(_2_6_io_y_sx),
    .io_y_sr(_2_6_io_y_sr),
    .io_y_pw(_2_6_io_y_pw),
    .io_y_px(_2_6_io_y_px),
    .io_y_pr(_2_6_io_y_pr),
    .io_y_pal(_2_6_io_y_pal),
    .io_y_paa(_2_6_io_y_paa),
    .io_y_eff(_2_6_io_y_eff),
    .io_y_c(_2_6_io_y_c)
  );
  _2_1 _2_7 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117713.4]
    .io_x_ppn(_2_7_io_x_ppn),
    .io_x_u(_2_7_io_x_u),
    .io_x_ae(_2_7_io_x_ae),
    .io_x_sw(_2_7_io_x_sw),
    .io_x_sx(_2_7_io_x_sx),
    .io_x_sr(_2_7_io_x_sr),
    .io_x_pw(_2_7_io_x_pw),
    .io_x_px(_2_7_io_x_px),
    .io_x_pr(_2_7_io_x_pr),
    .io_x_pal(_2_7_io_x_pal),
    .io_x_paa(_2_7_io_x_paa),
    .io_x_eff(_2_7_io_x_eff),
    .io_x_c(_2_7_io_x_c),
    .io_y_ppn(_2_7_io_y_ppn),
    .io_y_u(_2_7_io_y_u),
    .io_y_ae(_2_7_io_y_ae),
    .io_y_sw(_2_7_io_y_sw),
    .io_y_sx(_2_7_io_y_sx),
    .io_y_sr(_2_7_io_y_sr),
    .io_y_pw(_2_7_io_y_pw),
    .io_y_px(_2_7_io_y_px),
    .io_y_pr(_2_7_io_y_pr),
    .io_y_pal(_2_7_io_y_pal),
    .io_y_paa(_2_7_io_y_paa),
    .io_y_eff(_2_7_io_y_eff),
    .io_y_c(_2_7_io_y_c)
  );
  _2_1 _2_8 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117754.4]
    .io_x_ppn(_2_8_io_x_ppn),
    .io_x_u(_2_8_io_x_u),
    .io_x_ae(_2_8_io_x_ae),
    .io_x_sw(_2_8_io_x_sw),
    .io_x_sx(_2_8_io_x_sx),
    .io_x_sr(_2_8_io_x_sr),
    .io_x_pw(_2_8_io_x_pw),
    .io_x_px(_2_8_io_x_px),
    .io_x_pr(_2_8_io_x_pr),
    .io_x_pal(_2_8_io_x_pal),
    .io_x_paa(_2_8_io_x_paa),
    .io_x_eff(_2_8_io_x_eff),
    .io_x_c(_2_8_io_x_c),
    .io_y_ppn(_2_8_io_y_ppn),
    .io_y_u(_2_8_io_y_u),
    .io_y_ae(_2_8_io_y_ae),
    .io_y_sw(_2_8_io_y_sw),
    .io_y_sx(_2_8_io_y_sx),
    .io_y_sr(_2_8_io_y_sr),
    .io_y_pw(_2_8_io_y_pw),
    .io_y_px(_2_8_io_y_px),
    .io_y_pr(_2_8_io_y_pr),
    .io_y_pal(_2_8_io_y_pal),
    .io_y_paa(_2_8_io_y_paa),
    .io_y_eff(_2_8_io_y_eff),
    .io_y_c(_2_8_io_y_c)
  );
  _2_1 _2_9 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117794.4]
    .io_x_ppn(_2_9_io_x_ppn),
    .io_x_u(_2_9_io_x_u),
    .io_x_ae(_2_9_io_x_ae),
    .io_x_sw(_2_9_io_x_sw),
    .io_x_sx(_2_9_io_x_sx),
    .io_x_sr(_2_9_io_x_sr),
    .io_x_pw(_2_9_io_x_pw),
    .io_x_px(_2_9_io_x_px),
    .io_x_pr(_2_9_io_x_pr),
    .io_x_pal(_2_9_io_x_pal),
    .io_x_paa(_2_9_io_x_paa),
    .io_x_eff(_2_9_io_x_eff),
    .io_x_c(_2_9_io_x_c),
    .io_y_ppn(_2_9_io_y_ppn),
    .io_y_u(_2_9_io_y_u),
    .io_y_ae(_2_9_io_y_ae),
    .io_y_sw(_2_9_io_y_sw),
    .io_y_sx(_2_9_io_y_sx),
    .io_y_sr(_2_9_io_y_sr),
    .io_y_pw(_2_9_io_y_pw),
    .io_y_px(_2_9_io_y_px),
    .io_y_pr(_2_9_io_y_pr),
    .io_y_pal(_2_9_io_y_pal),
    .io_y_paa(_2_9_io_y_paa),
    .io_y_eff(_2_9_io_y_eff),
    .io_y_c(_2_9_io_y_c)
  );
  _2_1 _2_10 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117841.4]
    .io_x_ppn(_2_10_io_x_ppn),
    .io_x_u(_2_10_io_x_u),
    .io_x_ae(_2_10_io_x_ae),
    .io_x_sw(_2_10_io_x_sw),
    .io_x_sx(_2_10_io_x_sx),
    .io_x_sr(_2_10_io_x_sr),
    .io_x_pw(_2_10_io_x_pw),
    .io_x_px(_2_10_io_x_px),
    .io_x_pr(_2_10_io_x_pr),
    .io_x_pal(_2_10_io_x_pal),
    .io_x_paa(_2_10_io_x_paa),
    .io_x_eff(_2_10_io_x_eff),
    .io_x_c(_2_10_io_x_c),
    .io_y_ppn(_2_10_io_y_ppn),
    .io_y_u(_2_10_io_y_u),
    .io_y_ae(_2_10_io_y_ae),
    .io_y_sw(_2_10_io_y_sw),
    .io_y_sx(_2_10_io_y_sx),
    .io_y_sr(_2_10_io_y_sr),
    .io_y_pw(_2_10_io_y_pw),
    .io_y_px(_2_10_io_y_px),
    .io_y_pr(_2_10_io_y_pr),
    .io_y_pal(_2_10_io_y_pal),
    .io_y_paa(_2_10_io_y_paa),
    .io_y_eff(_2_10_io_y_eff),
    .io_y_c(_2_10_io_y_c)
  );
  _2_1 _2_11 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117888.4]
    .io_x_ppn(_2_11_io_x_ppn),
    .io_x_u(_2_11_io_x_u),
    .io_x_ae(_2_11_io_x_ae),
    .io_x_sw(_2_11_io_x_sw),
    .io_x_sx(_2_11_io_x_sx),
    .io_x_sr(_2_11_io_x_sr),
    .io_x_pw(_2_11_io_x_pw),
    .io_x_px(_2_11_io_x_px),
    .io_x_pr(_2_11_io_x_pr),
    .io_x_pal(_2_11_io_x_pal),
    .io_x_paa(_2_11_io_x_paa),
    .io_x_eff(_2_11_io_x_eff),
    .io_x_c(_2_11_io_x_c),
    .io_y_ppn(_2_11_io_y_ppn),
    .io_y_u(_2_11_io_y_u),
    .io_y_ae(_2_11_io_y_ae),
    .io_y_sw(_2_11_io_y_sw),
    .io_y_sx(_2_11_io_y_sx),
    .io_y_sr(_2_11_io_y_sr),
    .io_y_pw(_2_11_io_y_pw),
    .io_y_px(_2_11_io_y_px),
    .io_y_pr(_2_11_io_y_pr),
    .io_y_pal(_2_11_io_y_pal),
    .io_y_paa(_2_11_io_y_paa),
    .io_y_eff(_2_11_io_y_eff),
    .io_y_c(_2_11_io_y_c)
  );
  _2_1 _2_12 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117935.4]
    .io_x_ppn(_2_12_io_x_ppn),
    .io_x_u(_2_12_io_x_u),
    .io_x_ae(_2_12_io_x_ae),
    .io_x_sw(_2_12_io_x_sw),
    .io_x_sx(_2_12_io_x_sx),
    .io_x_sr(_2_12_io_x_sr),
    .io_x_pw(_2_12_io_x_pw),
    .io_x_px(_2_12_io_x_px),
    .io_x_pr(_2_12_io_x_pr),
    .io_x_pal(_2_12_io_x_pal),
    .io_x_paa(_2_12_io_x_paa),
    .io_x_eff(_2_12_io_x_eff),
    .io_x_c(_2_12_io_x_c),
    .io_y_ppn(_2_12_io_y_ppn),
    .io_y_u(_2_12_io_y_u),
    .io_y_ae(_2_12_io_y_ae),
    .io_y_sw(_2_12_io_y_sw),
    .io_y_sx(_2_12_io_y_sx),
    .io_y_sr(_2_12_io_y_sr),
    .io_y_pw(_2_12_io_y_pw),
    .io_y_px(_2_12_io_y_px),
    .io_y_pr(_2_12_io_y_pr),
    .io_y_pal(_2_12_io_y_pal),
    .io_y_paa(_2_12_io_y_paa),
    .io_y_eff(_2_12_io_y_eff),
    .io_y_c(_2_12_io_y_c)
  );
  _2_1 _2_13 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@117982.4]
    .io_x_ppn(_2_13_io_x_ppn),
    .io_x_u(_2_13_io_x_u),
    .io_x_ae(_2_13_io_x_ae),
    .io_x_sw(_2_13_io_x_sw),
    .io_x_sx(_2_13_io_x_sx),
    .io_x_sr(_2_13_io_x_sr),
    .io_x_pw(_2_13_io_x_pw),
    .io_x_px(_2_13_io_x_px),
    .io_x_pr(_2_13_io_x_pr),
    .io_x_pal(_2_13_io_x_pal),
    .io_x_paa(_2_13_io_x_paa),
    .io_x_eff(_2_13_io_x_eff),
    .io_x_c(_2_13_io_x_c),
    .io_y_ppn(_2_13_io_y_ppn),
    .io_y_u(_2_13_io_y_u),
    .io_y_ae(_2_13_io_y_ae),
    .io_y_sw(_2_13_io_y_sw),
    .io_y_sx(_2_13_io_y_sx),
    .io_y_sr(_2_13_io_y_sr),
    .io_y_pw(_2_13_io_y_pw),
    .io_y_px(_2_13_io_y_px),
    .io_y_pr(_2_13_io_y_pr),
    .io_y_pal(_2_13_io_y_pal),
    .io_y_paa(_2_13_io_y_paa),
    .io_y_eff(_2_13_io_y_eff),
    .io_y_c(_2_13_io_y_c)
  );
  _2_1 _2_14 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118447.4]
    .io_x_ppn(_2_14_io_x_ppn),
    .io_x_u(_2_14_io_x_u),
    .io_x_ae(_2_14_io_x_ae),
    .io_x_sw(_2_14_io_x_sw),
    .io_x_sx(_2_14_io_x_sx),
    .io_x_sr(_2_14_io_x_sr),
    .io_x_pw(_2_14_io_x_pw),
    .io_x_px(_2_14_io_x_px),
    .io_x_pr(_2_14_io_x_pr),
    .io_x_pal(_2_14_io_x_pal),
    .io_x_paa(_2_14_io_x_paa),
    .io_x_eff(_2_14_io_x_eff),
    .io_x_c(_2_14_io_x_c),
    .io_y_ppn(_2_14_io_y_ppn),
    .io_y_u(_2_14_io_y_u),
    .io_y_ae(_2_14_io_y_ae),
    .io_y_sw(_2_14_io_y_sw),
    .io_y_sx(_2_14_io_y_sx),
    .io_y_sr(_2_14_io_y_sr),
    .io_y_pw(_2_14_io_y_pw),
    .io_y_px(_2_14_io_y_px),
    .io_y_pr(_2_14_io_y_pr),
    .io_y_pal(_2_14_io_y_pal),
    .io_y_paa(_2_14_io_y_paa),
    .io_y_eff(_2_14_io_y_eff),
    .io_y_c(_2_14_io_y_c)
  );
  _2_1 _2_15 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118488.4]
    .io_x_ppn(_2_15_io_x_ppn),
    .io_x_u(_2_15_io_x_u),
    .io_x_ae(_2_15_io_x_ae),
    .io_x_sw(_2_15_io_x_sw),
    .io_x_sx(_2_15_io_x_sx),
    .io_x_sr(_2_15_io_x_sr),
    .io_x_pw(_2_15_io_x_pw),
    .io_x_px(_2_15_io_x_px),
    .io_x_pr(_2_15_io_x_pr),
    .io_x_pal(_2_15_io_x_pal),
    .io_x_paa(_2_15_io_x_paa),
    .io_x_eff(_2_15_io_x_eff),
    .io_x_c(_2_15_io_x_c),
    .io_y_ppn(_2_15_io_y_ppn),
    .io_y_u(_2_15_io_y_u),
    .io_y_ae(_2_15_io_y_ae),
    .io_y_sw(_2_15_io_y_sw),
    .io_y_sx(_2_15_io_y_sx),
    .io_y_sr(_2_15_io_y_sr),
    .io_y_pw(_2_15_io_y_pw),
    .io_y_px(_2_15_io_y_px),
    .io_y_pr(_2_15_io_y_pr),
    .io_y_pal(_2_15_io_y_pal),
    .io_y_paa(_2_15_io_y_paa),
    .io_y_eff(_2_15_io_y_eff),
    .io_y_c(_2_15_io_y_c)
  );
  _2_1 _2_16 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118529.4]
    .io_x_ppn(_2_16_io_x_ppn),
    .io_x_u(_2_16_io_x_u),
    .io_x_ae(_2_16_io_x_ae),
    .io_x_sw(_2_16_io_x_sw),
    .io_x_sx(_2_16_io_x_sx),
    .io_x_sr(_2_16_io_x_sr),
    .io_x_pw(_2_16_io_x_pw),
    .io_x_px(_2_16_io_x_px),
    .io_x_pr(_2_16_io_x_pr),
    .io_x_pal(_2_16_io_x_pal),
    .io_x_paa(_2_16_io_x_paa),
    .io_x_eff(_2_16_io_x_eff),
    .io_x_c(_2_16_io_x_c),
    .io_y_ppn(_2_16_io_y_ppn),
    .io_y_u(_2_16_io_y_u),
    .io_y_ae(_2_16_io_y_ae),
    .io_y_sw(_2_16_io_y_sw),
    .io_y_sx(_2_16_io_y_sx),
    .io_y_sr(_2_16_io_y_sr),
    .io_y_pw(_2_16_io_y_pw),
    .io_y_px(_2_16_io_y_px),
    .io_y_pr(_2_16_io_y_pr),
    .io_y_pal(_2_16_io_y_pal),
    .io_y_paa(_2_16_io_y_paa),
    .io_y_eff(_2_16_io_y_eff),
    .io_y_c(_2_16_io_y_c)
  );
  _2_1 _2_17 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118570.4]
    .io_x_ppn(_2_17_io_x_ppn),
    .io_x_u(_2_17_io_x_u),
    .io_x_ae(_2_17_io_x_ae),
    .io_x_sw(_2_17_io_x_sw),
    .io_x_sx(_2_17_io_x_sx),
    .io_x_sr(_2_17_io_x_sr),
    .io_x_pw(_2_17_io_x_pw),
    .io_x_px(_2_17_io_x_px),
    .io_x_pr(_2_17_io_x_pr),
    .io_x_pal(_2_17_io_x_pal),
    .io_x_paa(_2_17_io_x_paa),
    .io_x_eff(_2_17_io_x_eff),
    .io_x_c(_2_17_io_x_c),
    .io_y_ppn(_2_17_io_y_ppn),
    .io_y_u(_2_17_io_y_u),
    .io_y_ae(_2_17_io_y_ae),
    .io_y_sw(_2_17_io_y_sw),
    .io_y_sx(_2_17_io_y_sx),
    .io_y_sr(_2_17_io_y_sr),
    .io_y_pw(_2_17_io_y_pw),
    .io_y_px(_2_17_io_y_px),
    .io_y_pr(_2_17_io_y_pr),
    .io_y_pal(_2_17_io_y_pal),
    .io_y_paa(_2_17_io_y_paa),
    .io_y_eff(_2_17_io_y_eff),
    .io_y_c(_2_17_io_y_c)
  );
  _2_1 _2_18 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118611.4]
    .io_x_ppn(_2_18_io_x_ppn),
    .io_x_u(_2_18_io_x_u),
    .io_x_ae(_2_18_io_x_ae),
    .io_x_sw(_2_18_io_x_sw),
    .io_x_sx(_2_18_io_x_sx),
    .io_x_sr(_2_18_io_x_sr),
    .io_x_pw(_2_18_io_x_pw),
    .io_x_px(_2_18_io_x_px),
    .io_x_pr(_2_18_io_x_pr),
    .io_x_pal(_2_18_io_x_pal),
    .io_x_paa(_2_18_io_x_paa),
    .io_x_eff(_2_18_io_x_eff),
    .io_x_c(_2_18_io_x_c),
    .io_y_ppn(_2_18_io_y_ppn),
    .io_y_u(_2_18_io_y_u),
    .io_y_ae(_2_18_io_y_ae),
    .io_y_sw(_2_18_io_y_sw),
    .io_y_sx(_2_18_io_y_sx),
    .io_y_sr(_2_18_io_y_sr),
    .io_y_pw(_2_18_io_y_pw),
    .io_y_px(_2_18_io_y_px),
    .io_y_pr(_2_18_io_y_pr),
    .io_y_pal(_2_18_io_y_pal),
    .io_y_paa(_2_18_io_y_paa),
    .io_y_eff(_2_18_io_y_eff),
    .io_y_c(_2_18_io_y_c)
  );
  _2_1 _2_19 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118652.4]
    .io_x_ppn(_2_19_io_x_ppn),
    .io_x_u(_2_19_io_x_u),
    .io_x_ae(_2_19_io_x_ae),
    .io_x_sw(_2_19_io_x_sw),
    .io_x_sx(_2_19_io_x_sx),
    .io_x_sr(_2_19_io_x_sr),
    .io_x_pw(_2_19_io_x_pw),
    .io_x_px(_2_19_io_x_px),
    .io_x_pr(_2_19_io_x_pr),
    .io_x_pal(_2_19_io_x_pal),
    .io_x_paa(_2_19_io_x_paa),
    .io_x_eff(_2_19_io_x_eff),
    .io_x_c(_2_19_io_x_c),
    .io_y_ppn(_2_19_io_y_ppn),
    .io_y_u(_2_19_io_y_u),
    .io_y_ae(_2_19_io_y_ae),
    .io_y_sw(_2_19_io_y_sw),
    .io_y_sx(_2_19_io_y_sx),
    .io_y_sr(_2_19_io_y_sr),
    .io_y_pw(_2_19_io_y_pw),
    .io_y_px(_2_19_io_y_px),
    .io_y_pr(_2_19_io_y_pr),
    .io_y_pal(_2_19_io_y_pal),
    .io_y_paa(_2_19_io_y_paa),
    .io_y_eff(_2_19_io_y_eff),
    .io_y_c(_2_19_io_y_c)
  );
  _2_1 _2_20 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118693.4]
    .io_x_ppn(_2_20_io_x_ppn),
    .io_x_u(_2_20_io_x_u),
    .io_x_ae(_2_20_io_x_ae),
    .io_x_sw(_2_20_io_x_sw),
    .io_x_sx(_2_20_io_x_sx),
    .io_x_sr(_2_20_io_x_sr),
    .io_x_pw(_2_20_io_x_pw),
    .io_x_px(_2_20_io_x_px),
    .io_x_pr(_2_20_io_x_pr),
    .io_x_pal(_2_20_io_x_pal),
    .io_x_paa(_2_20_io_x_paa),
    .io_x_eff(_2_20_io_x_eff),
    .io_x_c(_2_20_io_x_c),
    .io_y_ppn(_2_20_io_y_ppn),
    .io_y_u(_2_20_io_y_u),
    .io_y_ae(_2_20_io_y_ae),
    .io_y_sw(_2_20_io_y_sw),
    .io_y_sx(_2_20_io_y_sx),
    .io_y_sr(_2_20_io_y_sr),
    .io_y_pw(_2_20_io_y_pw),
    .io_y_px(_2_20_io_y_px),
    .io_y_pr(_2_20_io_y_pr),
    .io_y_pal(_2_20_io_y_pal),
    .io_y_paa(_2_20_io_y_paa),
    .io_y_eff(_2_20_io_y_eff),
    .io_y_c(_2_20_io_y_c)
  );
  _2_1 _2_21 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118734.4]
    .io_x_ppn(_2_21_io_x_ppn),
    .io_x_u(_2_21_io_x_u),
    .io_x_ae(_2_21_io_x_ae),
    .io_x_sw(_2_21_io_x_sw),
    .io_x_sx(_2_21_io_x_sx),
    .io_x_sr(_2_21_io_x_sr),
    .io_x_pw(_2_21_io_x_pw),
    .io_x_px(_2_21_io_x_px),
    .io_x_pr(_2_21_io_x_pr),
    .io_x_pal(_2_21_io_x_pal),
    .io_x_paa(_2_21_io_x_paa),
    .io_x_eff(_2_21_io_x_eff),
    .io_x_c(_2_21_io_x_c),
    .io_y_ppn(_2_21_io_y_ppn),
    .io_y_u(_2_21_io_y_u),
    .io_y_ae(_2_21_io_y_ae),
    .io_y_sw(_2_21_io_y_sw),
    .io_y_sx(_2_21_io_y_sx),
    .io_y_sr(_2_21_io_y_sr),
    .io_y_pw(_2_21_io_y_pw),
    .io_y_px(_2_21_io_y_px),
    .io_y_pr(_2_21_io_y_pr),
    .io_y_pal(_2_21_io_y_pal),
    .io_y_paa(_2_21_io_y_paa),
    .io_y_eff(_2_21_io_y_eff),
    .io_y_c(_2_21_io_y_c)
  );
  _2_1 _2_22 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118774.4]
    .io_x_ppn(_2_22_io_x_ppn),
    .io_x_u(_2_22_io_x_u),
    .io_x_ae(_2_22_io_x_ae),
    .io_x_sw(_2_22_io_x_sw),
    .io_x_sx(_2_22_io_x_sx),
    .io_x_sr(_2_22_io_x_sr),
    .io_x_pw(_2_22_io_x_pw),
    .io_x_px(_2_22_io_x_px),
    .io_x_pr(_2_22_io_x_pr),
    .io_x_pal(_2_22_io_x_pal),
    .io_x_paa(_2_22_io_x_paa),
    .io_x_eff(_2_22_io_x_eff),
    .io_x_c(_2_22_io_x_c),
    .io_y_ppn(_2_22_io_y_ppn),
    .io_y_u(_2_22_io_y_u),
    .io_y_ae(_2_22_io_y_ae),
    .io_y_sw(_2_22_io_y_sw),
    .io_y_sx(_2_22_io_y_sx),
    .io_y_sr(_2_22_io_y_sr),
    .io_y_pw(_2_22_io_y_pw),
    .io_y_px(_2_22_io_y_px),
    .io_y_pr(_2_22_io_y_pr),
    .io_y_pal(_2_22_io_y_pal),
    .io_y_paa(_2_22_io_y_paa),
    .io_y_eff(_2_22_io_y_eff),
    .io_y_c(_2_22_io_y_c)
  );
  _2_1 _2_23 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118814.4]
    .io_x_ppn(_2_23_io_x_ppn),
    .io_x_u(_2_23_io_x_u),
    .io_x_ae(_2_23_io_x_ae),
    .io_x_sw(_2_23_io_x_sw),
    .io_x_sx(_2_23_io_x_sx),
    .io_x_sr(_2_23_io_x_sr),
    .io_x_pw(_2_23_io_x_pw),
    .io_x_px(_2_23_io_x_px),
    .io_x_pr(_2_23_io_x_pr),
    .io_x_pal(_2_23_io_x_pal),
    .io_x_paa(_2_23_io_x_paa),
    .io_x_eff(_2_23_io_x_eff),
    .io_x_c(_2_23_io_x_c),
    .io_y_ppn(_2_23_io_y_ppn),
    .io_y_u(_2_23_io_y_u),
    .io_y_ae(_2_23_io_y_ae),
    .io_y_sw(_2_23_io_y_sw),
    .io_y_sx(_2_23_io_y_sx),
    .io_y_sr(_2_23_io_y_sr),
    .io_y_pw(_2_23_io_y_pw),
    .io_y_px(_2_23_io_y_px),
    .io_y_pr(_2_23_io_y_pr),
    .io_y_pal(_2_23_io_y_pal),
    .io_y_paa(_2_23_io_y_paa),
    .io_y_eff(_2_23_io_y_eff),
    .io_y_c(_2_23_io_y_c)
  );
  _2_1 _2_24 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118854.4]
    .io_x_ppn(_2_24_io_x_ppn),
    .io_x_u(_2_24_io_x_u),
    .io_x_ae(_2_24_io_x_ae),
    .io_x_sw(_2_24_io_x_sw),
    .io_x_sx(_2_24_io_x_sx),
    .io_x_sr(_2_24_io_x_sr),
    .io_x_pw(_2_24_io_x_pw),
    .io_x_px(_2_24_io_x_px),
    .io_x_pr(_2_24_io_x_pr),
    .io_x_pal(_2_24_io_x_pal),
    .io_x_paa(_2_24_io_x_paa),
    .io_x_eff(_2_24_io_x_eff),
    .io_x_c(_2_24_io_x_c),
    .io_y_ppn(_2_24_io_y_ppn),
    .io_y_u(_2_24_io_y_u),
    .io_y_ae(_2_24_io_y_ae),
    .io_y_sw(_2_24_io_y_sw),
    .io_y_sx(_2_24_io_y_sx),
    .io_y_sr(_2_24_io_y_sr),
    .io_y_pw(_2_24_io_y_pw),
    .io_y_px(_2_24_io_y_px),
    .io_y_pr(_2_24_io_y_pr),
    .io_y_pal(_2_24_io_y_pal),
    .io_y_paa(_2_24_io_y_paa),
    .io_y_eff(_2_24_io_y_eff),
    .io_y_c(_2_24_io_y_c)
  );
  _2_1 _2_25 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118894.4]
    .io_x_ppn(_2_25_io_x_ppn),
    .io_x_u(_2_25_io_x_u),
    .io_x_ae(_2_25_io_x_ae),
    .io_x_sw(_2_25_io_x_sw),
    .io_x_sx(_2_25_io_x_sx),
    .io_x_sr(_2_25_io_x_sr),
    .io_x_pw(_2_25_io_x_pw),
    .io_x_px(_2_25_io_x_px),
    .io_x_pr(_2_25_io_x_pr),
    .io_x_pal(_2_25_io_x_pal),
    .io_x_paa(_2_25_io_x_paa),
    .io_x_eff(_2_25_io_x_eff),
    .io_x_c(_2_25_io_x_c),
    .io_y_ppn(_2_25_io_y_ppn),
    .io_y_u(_2_25_io_y_u),
    .io_y_ae(_2_25_io_y_ae),
    .io_y_sw(_2_25_io_y_sw),
    .io_y_sx(_2_25_io_y_sx),
    .io_y_sr(_2_25_io_y_sr),
    .io_y_pw(_2_25_io_y_pw),
    .io_y_px(_2_25_io_y_px),
    .io_y_pr(_2_25_io_y_pr),
    .io_y_pal(_2_25_io_y_pal),
    .io_y_paa(_2_25_io_y_paa),
    .io_y_eff(_2_25_io_y_eff),
    .io_y_c(_2_25_io_y_c)
  );
  _2_1 _2_26 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118934.4]
    .io_x_ppn(_2_26_io_x_ppn),
    .io_x_u(_2_26_io_x_u),
    .io_x_ae(_2_26_io_x_ae),
    .io_x_sw(_2_26_io_x_sw),
    .io_x_sx(_2_26_io_x_sx),
    .io_x_sr(_2_26_io_x_sr),
    .io_x_pw(_2_26_io_x_pw),
    .io_x_px(_2_26_io_x_px),
    .io_x_pr(_2_26_io_x_pr),
    .io_x_pal(_2_26_io_x_pal),
    .io_x_paa(_2_26_io_x_paa),
    .io_x_eff(_2_26_io_x_eff),
    .io_x_c(_2_26_io_x_c),
    .io_y_ppn(_2_26_io_y_ppn),
    .io_y_u(_2_26_io_y_u),
    .io_y_ae(_2_26_io_y_ae),
    .io_y_sw(_2_26_io_y_sw),
    .io_y_sx(_2_26_io_y_sx),
    .io_y_sr(_2_26_io_y_sr),
    .io_y_pw(_2_26_io_y_pw),
    .io_y_px(_2_26_io_y_px),
    .io_y_pr(_2_26_io_y_pr),
    .io_y_pal(_2_26_io_y_pal),
    .io_y_paa(_2_26_io_y_paa),
    .io_y_eff(_2_26_io_y_eff),
    .io_y_c(_2_26_io_y_c)
  );
  _2_1 _2_27 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@118975.4]
    .io_x_ppn(_2_27_io_x_ppn),
    .io_x_u(_2_27_io_x_u),
    .io_x_ae(_2_27_io_x_ae),
    .io_x_sw(_2_27_io_x_sw),
    .io_x_sx(_2_27_io_x_sx),
    .io_x_sr(_2_27_io_x_sr),
    .io_x_pw(_2_27_io_x_pw),
    .io_x_px(_2_27_io_x_px),
    .io_x_pr(_2_27_io_x_pr),
    .io_x_pal(_2_27_io_x_pal),
    .io_x_paa(_2_27_io_x_paa),
    .io_x_eff(_2_27_io_x_eff),
    .io_x_c(_2_27_io_x_c),
    .io_y_ppn(_2_27_io_y_ppn),
    .io_y_u(_2_27_io_y_u),
    .io_y_ae(_2_27_io_y_ae),
    .io_y_sw(_2_27_io_y_sw),
    .io_y_sx(_2_27_io_y_sx),
    .io_y_sr(_2_27_io_y_sr),
    .io_y_pw(_2_27_io_y_pw),
    .io_y_px(_2_27_io_y_px),
    .io_y_pr(_2_27_io_y_pr),
    .io_y_pal(_2_27_io_y_pal),
    .io_y_paa(_2_27_io_y_paa),
    .io_y_eff(_2_27_io_y_eff),
    .io_y_c(_2_27_io_y_c)
  );
  _2_1 _2_28 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119016.4]
    .io_x_ppn(_2_28_io_x_ppn),
    .io_x_u(_2_28_io_x_u),
    .io_x_ae(_2_28_io_x_ae),
    .io_x_sw(_2_28_io_x_sw),
    .io_x_sx(_2_28_io_x_sx),
    .io_x_sr(_2_28_io_x_sr),
    .io_x_pw(_2_28_io_x_pw),
    .io_x_px(_2_28_io_x_px),
    .io_x_pr(_2_28_io_x_pr),
    .io_x_pal(_2_28_io_x_pal),
    .io_x_paa(_2_28_io_x_paa),
    .io_x_eff(_2_28_io_x_eff),
    .io_x_c(_2_28_io_x_c),
    .io_y_ppn(_2_28_io_y_ppn),
    .io_y_u(_2_28_io_y_u),
    .io_y_ae(_2_28_io_y_ae),
    .io_y_sw(_2_28_io_y_sw),
    .io_y_sx(_2_28_io_y_sx),
    .io_y_sr(_2_28_io_y_sr),
    .io_y_pw(_2_28_io_y_pw),
    .io_y_px(_2_28_io_y_px),
    .io_y_pr(_2_28_io_y_pr),
    .io_y_pal(_2_28_io_y_pal),
    .io_y_paa(_2_28_io_y_paa),
    .io_y_eff(_2_28_io_y_eff),
    .io_y_c(_2_28_io_y_c)
  );
  _2_1 _2_29 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119057.4]
    .io_x_ppn(_2_29_io_x_ppn),
    .io_x_u(_2_29_io_x_u),
    .io_x_ae(_2_29_io_x_ae),
    .io_x_sw(_2_29_io_x_sw),
    .io_x_sx(_2_29_io_x_sx),
    .io_x_sr(_2_29_io_x_sr),
    .io_x_pw(_2_29_io_x_pw),
    .io_x_px(_2_29_io_x_px),
    .io_x_pr(_2_29_io_x_pr),
    .io_x_pal(_2_29_io_x_pal),
    .io_x_paa(_2_29_io_x_paa),
    .io_x_eff(_2_29_io_x_eff),
    .io_x_c(_2_29_io_x_c),
    .io_y_ppn(_2_29_io_y_ppn),
    .io_y_u(_2_29_io_y_u),
    .io_y_ae(_2_29_io_y_ae),
    .io_y_sw(_2_29_io_y_sw),
    .io_y_sx(_2_29_io_y_sx),
    .io_y_sr(_2_29_io_y_sr),
    .io_y_pw(_2_29_io_y_pw),
    .io_y_px(_2_29_io_y_px),
    .io_y_pr(_2_29_io_y_pr),
    .io_y_pal(_2_29_io_y_pal),
    .io_y_paa(_2_29_io_y_paa),
    .io_y_eff(_2_29_io_y_eff),
    .io_y_c(_2_29_io_y_c)
  );
  _2_1 _2_30 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119098.4]
    .io_x_ppn(_2_30_io_x_ppn),
    .io_x_u(_2_30_io_x_u),
    .io_x_ae(_2_30_io_x_ae),
    .io_x_sw(_2_30_io_x_sw),
    .io_x_sx(_2_30_io_x_sx),
    .io_x_sr(_2_30_io_x_sr),
    .io_x_pw(_2_30_io_x_pw),
    .io_x_px(_2_30_io_x_px),
    .io_x_pr(_2_30_io_x_pr),
    .io_x_pal(_2_30_io_x_pal),
    .io_x_paa(_2_30_io_x_paa),
    .io_x_eff(_2_30_io_x_eff),
    .io_x_c(_2_30_io_x_c),
    .io_y_ppn(_2_30_io_y_ppn),
    .io_y_u(_2_30_io_y_u),
    .io_y_ae(_2_30_io_y_ae),
    .io_y_sw(_2_30_io_y_sw),
    .io_y_sx(_2_30_io_y_sx),
    .io_y_sr(_2_30_io_y_sr),
    .io_y_pw(_2_30_io_y_pw),
    .io_y_px(_2_30_io_y_px),
    .io_y_pr(_2_30_io_y_pr),
    .io_y_pal(_2_30_io_y_pal),
    .io_y_paa(_2_30_io_y_paa),
    .io_y_eff(_2_30_io_y_eff),
    .io_y_c(_2_30_io_y_c)
  );
  _2_1 _2_31 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119139.4]
    .io_x_ppn(_2_31_io_x_ppn),
    .io_x_u(_2_31_io_x_u),
    .io_x_ae(_2_31_io_x_ae),
    .io_x_sw(_2_31_io_x_sw),
    .io_x_sx(_2_31_io_x_sx),
    .io_x_sr(_2_31_io_x_sr),
    .io_x_pw(_2_31_io_x_pw),
    .io_x_px(_2_31_io_x_px),
    .io_x_pr(_2_31_io_x_pr),
    .io_x_pal(_2_31_io_x_pal),
    .io_x_paa(_2_31_io_x_paa),
    .io_x_eff(_2_31_io_x_eff),
    .io_x_c(_2_31_io_x_c),
    .io_y_ppn(_2_31_io_y_ppn),
    .io_y_u(_2_31_io_y_u),
    .io_y_ae(_2_31_io_y_ae),
    .io_y_sw(_2_31_io_y_sw),
    .io_y_sx(_2_31_io_y_sx),
    .io_y_sr(_2_31_io_y_sr),
    .io_y_pw(_2_31_io_y_pw),
    .io_y_px(_2_31_io_y_px),
    .io_y_pr(_2_31_io_y_pr),
    .io_y_pal(_2_31_io_y_pal),
    .io_y_paa(_2_31_io_y_paa),
    .io_y_eff(_2_31_io_y_eff),
    .io_y_c(_2_31_io_y_c)
  );
  _2_1 _2_32 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119180.4]
    .io_x_ppn(_2_32_io_x_ppn),
    .io_x_u(_2_32_io_x_u),
    .io_x_ae(_2_32_io_x_ae),
    .io_x_sw(_2_32_io_x_sw),
    .io_x_sx(_2_32_io_x_sx),
    .io_x_sr(_2_32_io_x_sr),
    .io_x_pw(_2_32_io_x_pw),
    .io_x_px(_2_32_io_x_px),
    .io_x_pr(_2_32_io_x_pr),
    .io_x_pal(_2_32_io_x_pal),
    .io_x_paa(_2_32_io_x_paa),
    .io_x_eff(_2_32_io_x_eff),
    .io_x_c(_2_32_io_x_c),
    .io_y_ppn(_2_32_io_y_ppn),
    .io_y_u(_2_32_io_y_u),
    .io_y_ae(_2_32_io_y_ae),
    .io_y_sw(_2_32_io_y_sw),
    .io_y_sx(_2_32_io_y_sx),
    .io_y_sr(_2_32_io_y_sr),
    .io_y_pw(_2_32_io_y_pw),
    .io_y_px(_2_32_io_y_px),
    .io_y_pr(_2_32_io_y_pr),
    .io_y_pal(_2_32_io_y_pal),
    .io_y_paa(_2_32_io_y_paa),
    .io_y_eff(_2_32_io_y_eff),
    .io_y_c(_2_32_io_y_c)
  );
  _2_1 _2_33 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119221.4]
    .io_x_ppn(_2_33_io_x_ppn),
    .io_x_u(_2_33_io_x_u),
    .io_x_ae(_2_33_io_x_ae),
    .io_x_sw(_2_33_io_x_sw),
    .io_x_sx(_2_33_io_x_sx),
    .io_x_sr(_2_33_io_x_sr),
    .io_x_pw(_2_33_io_x_pw),
    .io_x_px(_2_33_io_x_px),
    .io_x_pr(_2_33_io_x_pr),
    .io_x_pal(_2_33_io_x_pal),
    .io_x_paa(_2_33_io_x_paa),
    .io_x_eff(_2_33_io_x_eff),
    .io_x_c(_2_33_io_x_c),
    .io_y_ppn(_2_33_io_y_ppn),
    .io_y_u(_2_33_io_y_u),
    .io_y_ae(_2_33_io_y_ae),
    .io_y_sw(_2_33_io_y_sw),
    .io_y_sx(_2_33_io_y_sx),
    .io_y_sr(_2_33_io_y_sr),
    .io_y_pw(_2_33_io_y_pw),
    .io_y_px(_2_33_io_y_px),
    .io_y_pr(_2_33_io_y_pr),
    .io_y_pal(_2_33_io_y_pal),
    .io_y_paa(_2_33_io_y_paa),
    .io_y_eff(_2_33_io_y_eff),
    .io_y_c(_2_33_io_y_c)
  );
  _2_1 _2_34 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119262.4]
    .io_x_ppn(_2_34_io_x_ppn),
    .io_x_u(_2_34_io_x_u),
    .io_x_ae(_2_34_io_x_ae),
    .io_x_sw(_2_34_io_x_sw),
    .io_x_sx(_2_34_io_x_sx),
    .io_x_sr(_2_34_io_x_sr),
    .io_x_pw(_2_34_io_x_pw),
    .io_x_px(_2_34_io_x_px),
    .io_x_pr(_2_34_io_x_pr),
    .io_x_pal(_2_34_io_x_pal),
    .io_x_paa(_2_34_io_x_paa),
    .io_x_eff(_2_34_io_x_eff),
    .io_x_c(_2_34_io_x_c),
    .io_y_ppn(_2_34_io_y_ppn),
    .io_y_u(_2_34_io_y_u),
    .io_y_ae(_2_34_io_y_ae),
    .io_y_sw(_2_34_io_y_sw),
    .io_y_sx(_2_34_io_y_sx),
    .io_y_sr(_2_34_io_y_sr),
    .io_y_pw(_2_34_io_y_pw),
    .io_y_px(_2_34_io_y_px),
    .io_y_pr(_2_34_io_y_pr),
    .io_y_pal(_2_34_io_y_pal),
    .io_y_paa(_2_34_io_y_paa),
    .io_y_eff(_2_34_io_y_eff),
    .io_y_c(_2_34_io_y_c)
  );
  _2_1 _2_35 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119302.4]
    .io_x_ppn(_2_35_io_x_ppn),
    .io_x_u(_2_35_io_x_u),
    .io_x_ae(_2_35_io_x_ae),
    .io_x_sw(_2_35_io_x_sw),
    .io_x_sx(_2_35_io_x_sx),
    .io_x_sr(_2_35_io_x_sr),
    .io_x_pw(_2_35_io_x_pw),
    .io_x_px(_2_35_io_x_px),
    .io_x_pr(_2_35_io_x_pr),
    .io_x_pal(_2_35_io_x_pal),
    .io_x_paa(_2_35_io_x_paa),
    .io_x_eff(_2_35_io_x_eff),
    .io_x_c(_2_35_io_x_c),
    .io_y_ppn(_2_35_io_y_ppn),
    .io_y_u(_2_35_io_y_u),
    .io_y_ae(_2_35_io_y_ae),
    .io_y_sw(_2_35_io_y_sw),
    .io_y_sx(_2_35_io_y_sx),
    .io_y_sr(_2_35_io_y_sr),
    .io_y_pw(_2_35_io_y_pw),
    .io_y_px(_2_35_io_y_px),
    .io_y_pr(_2_35_io_y_pr),
    .io_y_pal(_2_35_io_y_pal),
    .io_y_paa(_2_35_io_y_paa),
    .io_y_eff(_2_35_io_y_eff),
    .io_y_c(_2_35_io_y_c)
  );
  _2_1 _2_36 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119342.4]
    .io_x_ppn(_2_36_io_x_ppn),
    .io_x_u(_2_36_io_x_u),
    .io_x_ae(_2_36_io_x_ae),
    .io_x_sw(_2_36_io_x_sw),
    .io_x_sx(_2_36_io_x_sx),
    .io_x_sr(_2_36_io_x_sr),
    .io_x_pw(_2_36_io_x_pw),
    .io_x_px(_2_36_io_x_px),
    .io_x_pr(_2_36_io_x_pr),
    .io_x_pal(_2_36_io_x_pal),
    .io_x_paa(_2_36_io_x_paa),
    .io_x_eff(_2_36_io_x_eff),
    .io_x_c(_2_36_io_x_c),
    .io_y_ppn(_2_36_io_y_ppn),
    .io_y_u(_2_36_io_y_u),
    .io_y_ae(_2_36_io_y_ae),
    .io_y_sw(_2_36_io_y_sw),
    .io_y_sx(_2_36_io_y_sx),
    .io_y_sr(_2_36_io_y_sr),
    .io_y_pw(_2_36_io_y_pw),
    .io_y_px(_2_36_io_y_px),
    .io_y_pr(_2_36_io_y_pr),
    .io_y_pal(_2_36_io_y_pal),
    .io_y_paa(_2_36_io_y_paa),
    .io_y_eff(_2_36_io_y_eff),
    .io_y_c(_2_36_io_y_c)
  );
  _2_1 _2_37 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119382.4]
    .io_x_ppn(_2_37_io_x_ppn),
    .io_x_u(_2_37_io_x_u),
    .io_x_ae(_2_37_io_x_ae),
    .io_x_sw(_2_37_io_x_sw),
    .io_x_sx(_2_37_io_x_sx),
    .io_x_sr(_2_37_io_x_sr),
    .io_x_pw(_2_37_io_x_pw),
    .io_x_px(_2_37_io_x_px),
    .io_x_pr(_2_37_io_x_pr),
    .io_x_pal(_2_37_io_x_pal),
    .io_x_paa(_2_37_io_x_paa),
    .io_x_eff(_2_37_io_x_eff),
    .io_x_c(_2_37_io_x_c),
    .io_y_ppn(_2_37_io_y_ppn),
    .io_y_u(_2_37_io_y_u),
    .io_y_ae(_2_37_io_y_ae),
    .io_y_sw(_2_37_io_y_sw),
    .io_y_sx(_2_37_io_y_sx),
    .io_y_sr(_2_37_io_y_sr),
    .io_y_pw(_2_37_io_y_pw),
    .io_y_px(_2_37_io_y_px),
    .io_y_pr(_2_37_io_y_pr),
    .io_y_pal(_2_37_io_y_pal),
    .io_y_paa(_2_37_io_y_paa),
    .io_y_eff(_2_37_io_y_eff),
    .io_y_c(_2_37_io_y_c)
  );
  _2_1 _2_38 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@119422.4]
    .io_x_ppn(_2_38_io_x_ppn),
    .io_x_u(_2_38_io_x_u),
    .io_x_ae(_2_38_io_x_ae),
    .io_x_sw(_2_38_io_x_sw),
    .io_x_sx(_2_38_io_x_sx),
    .io_x_sr(_2_38_io_x_sr),
    .io_x_pw(_2_38_io_x_pw),
    .io_x_px(_2_38_io_x_px),
    .io_x_pr(_2_38_io_x_pr),
    .io_x_pal(_2_38_io_x_pal),
    .io_x_paa(_2_38_io_x_paa),
    .io_x_eff(_2_38_io_x_eff),
    .io_x_c(_2_38_io_x_c),
    .io_y_ppn(_2_38_io_y_ppn),
    .io_y_u(_2_38_io_y_u),
    .io_y_ae(_2_38_io_y_ae),
    .io_y_sw(_2_38_io_y_sw),
    .io_y_sx(_2_38_io_y_sx),
    .io_y_sr(_2_38_io_y_sr),
    .io_y_pw(_2_38_io_y_pw),
    .io_y_px(_2_38_io_y_px),
    .io_y_pr(_2_38_io_y_pr),
    .io_y_pal(_2_38_io_y_pal),
    .io_y_paa(_2_38_io_y_paa),
    .io_y_eff(_2_38_io_y_eff),
    .io_y_c(_2_38_io_y_c)
  );
  assign priv_s = io_ptw_status_dprv[0]; // @[TLB.scala 176:20:freechips.rocketchip.system.DefaultRV32Config.fir@116732.4]
  assign priv_uses_vm = io_ptw_status_dprv <= 2'h1; // @[TLB.scala 177:27:freechips.rocketchip.system.DefaultRV32Config.fir@116733.4]
  assign _T_2 = io_ptw_ptbr_mode & priv_uses_vm; // @[TLB.scala 178:83:freechips.rocketchip.system.DefaultRV32Config.fir@116736.4]
  assign _T_3 = io_req_bits_passthrough == 1'h0; // @[TLB.scala 178:102:freechips.rocketchip.system.DefaultRV32Config.fir@116737.4]
  assign vm_enabled = _T_2 & _T_3; // @[TLB.scala 178:99:freechips.rocketchip.system.DefaultRV32Config.fir@116738.4]
  assign vpn = io_req_bits_vaddr[31:12]; // @[TLB.scala 181:30:freechips.rocketchip.system.DefaultRV32Config.fir@116739.4]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 182:44:freechips.rocketchip.system.DefaultRV32Config.fir@116740.4]
  assign _T_4 = state == 2'h1; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@116742.4]
  assign _T_5 = state == 2'h3; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@116743.4]
  assign invalidate_refill = _T_4 | _T_5; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@116744.4]
  assign _T_21 = special_entry_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@116775.4]
  assign _T_24 = _2_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@116786.4]
  assign _T_25 = special_entry_level < 1'h1; // @[TLB.scala 121:30:freechips.rocketchip.system.DefaultRV32Config.fir@116787.4]
  assign _T_27 = _T_25 ? vpn : 20'h0; // @[TLB.scala 122:30:freechips.rocketchip.system.DefaultRV32Config.fir@116789.4]
  assign _T_28 = _T_27 | _2_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@116790.4]
  assign _T_29 = _T_28[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@116791.4]
  assign _T_30 = {_T_24,_T_29}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@116792.4]
  assign _T_31 = io_req_bits_vaddr[31:12]; // @[TLB.scala 186:123:freechips.rocketchip.system.DefaultRV32Config.fir@116793.4]
  assign _T_32 = vm_enabled ? _T_30 : _T_31; // @[TLB.scala 186:20:freechips.rocketchip.system.DefaultRV32Config.fir@116794.4]
  assign mpu_ppn = io_ptw_resp_valid ? refill_ppn : _T_32; // @[TLB.scala 185:20:freechips.rocketchip.system.DefaultRV32Config.fir@116795.4]
  assign _T_33 = io_req_bits_vaddr[11:0]; // @[TLB.scala 187:52:freechips.rocketchip.system.DefaultRV32Config.fir@116796.4]
  assign mpu_physaddr = {mpu_ppn,_T_33}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@116797.4]
  assign _T_34 = io_ptw_resp_valid | io_req_bits_passthrough; // @[TLB.scala 188:56:freechips.rocketchip.system.DefaultRV32Config.fir@116798.4]
  assign _T_36 = {io_ptw_status_debug,io_ptw_status_dprv}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@116800.4]
  assign mpu_priv = _T_34 ? 3'h1 : _T_36; // @[TLB.scala 188:27:freechips.rocketchip.system.DefaultRV32Config.fir@116801.4]
  assign _T_37 = mpu_physaddr ^ 32'h3000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116817.4]
  assign _T_38 = {1'b0,$signed(_T_37)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116818.4]
  assign _T_39 = $signed(_T_38) & $signed(-33'sh1000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116819.4]
  assign _T_40 = $signed(_T_39); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116820.4]
  assign _T_41 = $signed(_T_40) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116821.4]
  assign _T_42 = mpu_physaddr ^ 32'hc000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116822.4]
  assign _T_43 = {1'b0,$signed(_T_42)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116823.4]
  assign _T_44 = $signed(_T_43) & $signed(-33'sh4000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116824.4]
  assign _T_45 = $signed(_T_44); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116825.4]
  assign _T_46 = $signed(_T_45) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116826.4]
  assign _T_47 = mpu_physaddr ^ 32'h2000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116827.4]
  assign _T_48 = {1'b0,$signed(_T_47)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116828.4]
  assign _T_49 = $signed(_T_48) & $signed(-33'sh10000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116829.4]
  assign _T_50 = $signed(_T_49); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116830.4]
  assign _T_51 = $signed(_T_50) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116831.4]
  assign _T_53 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116833.4]
  assign _T_54 = $signed(_T_53) & $signed(-33'sh1000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116834.4]
  assign _T_55 = $signed(_T_54); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116835.4]
  assign _T_56 = $signed(_T_55) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116836.4]
  assign _T_57 = mpu_physaddr ^ 32'h10000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116837.4]
  assign _T_58 = {1'b0,$signed(_T_57)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116838.4]
  assign _T_59 = $signed(_T_58) & $signed(-33'sh10000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116839.4]
  assign _T_60 = $signed(_T_59); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116840.4]
  assign _T_61 = $signed(_T_60) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116841.4]
  assign _T_62 = mpu_physaddr ^ 32'h80000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116842.4]
  assign _T_63 = {1'b0,$signed(_T_62)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116843.4]
  assign _T_64 = $signed(_T_63) & $signed(-33'sh10000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116844.4]
  assign _T_65 = $signed(_T_64); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116845.4]
  assign _T_66 = $signed(_T_65) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116846.4]
  assign _T_67 = mpu_physaddr ^ 32'h60000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116847.4]
  assign _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116848.4]
  assign _T_69 = $signed(_T_68) & $signed(-33'sh20000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116849.4]
  assign _T_70 = $signed(_T_69); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116850.4]
  assign _T_71 = $signed(_T_70) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116851.4]
  assign _T_73 = _T_41 | _T_46; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116861.4]
  assign _T_74 = _T_73 | _T_51; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116862.4]
  assign _T_75 = _T_74 | _T_56; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116863.4]
  assign _T_76 = _T_75 | _T_61; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116864.4]
  assign _T_77 = _T_76 | _T_66; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116865.4]
  assign legal_address = _T_77 | _T_71; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@116866.4]
  assign _T_85 = $signed(_T_63) & $signed(33'sh80000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116874.4]
  assign _T_86 = $signed(_T_85); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116875.4]
  assign _T_87 = $signed(_T_86) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116876.4]
  assign cacheable = legal_address & _T_87; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@116882.4]
  assign _T_142 = mpu_physaddr ^ 32'h8000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@116934.4]
  assign _T_143 = {1'b0,$signed(_T_142)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@116935.4]
  assign _T_144 = $signed(_T_143) & $signed(33'shc8000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116936.4]
  assign _T_145 = $signed(_T_144); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116937.4]
  assign _T_146 = $signed(_T_145) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116938.4]
  assign _T_163 = $signed(_T_53) & $signed(33'shc8010000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116955.4]
  assign _T_164 = $signed(_T_163); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@116956.4]
  assign _T_165 = $signed(_T_164) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@116957.4]
  assign _T_172 = _T_165 | _T_146; // @[TLBPermissions.scala 82:66:freechips.rocketchip.system.DefaultRV32Config.fir@116964.4]
  assign _T_185 = mpu_priv <= 3'h3; // @[TLB.scala 199:39:freechips.rocketchip.system.DefaultRV32Config.fir@116977.4]
  assign deny_access_to_debug = _T_185 & _T_56; // @[TLB.scala 199:48:freechips.rocketchip.system.DefaultRV32Config.fir@116983.4]
  assign _T_197 = deny_access_to_debug == 1'h0; // @[TLB.scala 200:44:freechips.rocketchip.system.DefaultRV32Config.fir@116990.4]
  assign _T_198 = legal_address & _T_197; // @[TLB.scala 200:41:freechips.rocketchip.system.DefaultRV32Config.fir@116991.4]
  assign prot_r = _T_198 & pmp_io_r; // @[TLB.scala 200:66:freechips.rocketchip.system.DefaultRV32Config.fir@116992.4]
  assign _T_211 = $signed(_T_63) & $signed(33'shc0000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117005.4]
  assign _T_212 = $signed(_T_211); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117006.4]
  assign _T_213 = $signed(_T_212) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117007.4]
  assign _T_214 = mpu_physaddr ^ 32'h40000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@117008.4]
  assign _T_215 = {1'b0,$signed(_T_214)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@117009.4]
  assign _T_216 = $signed(_T_215) & $signed(33'shc0000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117010.4]
  assign _T_217 = $signed(_T_216); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117011.4]
  assign _T_218 = $signed(_T_217) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117012.4]
  assign _T_220 = _T_172 | _T_213; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117014.4]
  assign _T_221 = _T_220 | _T_218; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117015.4]
  assign _T_231 = legal_address & _T_221; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@117026.4]
  assign _T_233 = _T_231 & _T_197; // @[TLB.scala 201:45:freechips.rocketchip.system.DefaultRV32Config.fir@117028.4]
  assign prot_w = _T_233 & pmp_io_w; // @[TLB.scala 201:70:freechips.rocketchip.system.DefaultRV32Config.fir@117029.4]
  assign prot_al = legal_address & _T_172; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@117063.4]
  assign _T_300 = $signed(_T_53) & $signed(33'shca000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117100.4]
  assign _T_301 = $signed(_T_300); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117101.4]
  assign _T_302 = $signed(_T_301) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117102.4]
  assign _T_313 = _T_302 | _T_213; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117113.4]
  assign _T_314 = _T_313 | _T_218; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117114.4]
  assign _T_330 = legal_address & _T_314; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@117131.4]
  assign _T_332 = _T_330 & _T_197; // @[TLB.scala 204:40:freechips.rocketchip.system.DefaultRV32Config.fir@117133.4]
  assign prot_x = _T_332 & pmp_io_x; // @[TLB.scala 204:65:freechips.rocketchip.system.DefaultRV32Config.fir@117134.4]
  assign _T_357 = $signed(_T_48) & $signed(33'shca010000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117159.4]
  assign _T_358 = $signed(_T_357); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117160.4]
  assign _T_359 = $signed(_T_358) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117161.4]
  assign _T_362 = $signed(_T_53) & $signed(33'shca012000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117164.4]
  assign _T_363 = $signed(_T_362); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@117165.4]
  assign _T_364 = $signed(_T_363) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@117166.4]
  assign _T_370 = _T_146 | _T_359; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117172.4]
  assign _T_371 = _T_370 | _T_364; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117173.4]
  assign _T_372 = _T_371 | _T_218; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@117174.4]
  assign prot_eff = legal_address & _T_372; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@117180.4]
  assign _T_377 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117181.4]
  assign _T_378 = _T_377 | sectored_entries_0_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117182.4]
  assign _T_379 = _T_378 | sectored_entries_0_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117183.4]
  assign _T_380 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117184.4]
  assign _T_381 = _T_380[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117185.4]
  assign _T_382 = _T_381 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117186.4]
  assign sector_hits_0 = _T_379 & _T_382; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117187.4]
  assign _T_383 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117188.4]
  assign _T_384 = _T_383 | sectored_entries_1_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117189.4]
  assign _T_385 = _T_384 | sectored_entries_1_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117190.4]
  assign _T_386 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117191.4]
  assign _T_387 = _T_386[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117192.4]
  assign _T_388 = _T_387 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117193.4]
  assign sector_hits_1 = _T_385 & _T_388; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117194.4]
  assign _T_389 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117195.4]
  assign _T_390 = _T_389 | sectored_entries_2_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117196.4]
  assign _T_391 = _T_390 | sectored_entries_2_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117197.4]
  assign _T_392 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117198.4]
  assign _T_393 = _T_392[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117199.4]
  assign _T_394 = _T_393 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117200.4]
  assign sector_hits_2 = _T_391 & _T_394; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117201.4]
  assign _T_395 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117202.4]
  assign _T_396 = _T_395 | sectored_entries_3_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117203.4]
  assign _T_397 = _T_396 | sectored_entries_3_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117204.4]
  assign _T_398 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117205.4]
  assign _T_399 = _T_398[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117206.4]
  assign _T_400 = _T_399 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117207.4]
  assign sector_hits_3 = _T_397 & _T_400; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117208.4]
  assign _T_401 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117209.4]
  assign _T_402 = _T_401 | sectored_entries_4_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117210.4]
  assign _T_403 = _T_402 | sectored_entries_4_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117211.4]
  assign _T_404 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117212.4]
  assign _T_405 = _T_404[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117213.4]
  assign _T_406 = _T_405 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117214.4]
  assign sector_hits_4 = _T_403 & _T_406; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117215.4]
  assign _T_407 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117216.4]
  assign _T_408 = _T_407 | sectored_entries_5_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117217.4]
  assign _T_409 = _T_408 | sectored_entries_5_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117218.4]
  assign _T_410 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117219.4]
  assign _T_411 = _T_410[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117220.4]
  assign _T_412 = _T_411 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117221.4]
  assign sector_hits_5 = _T_409 & _T_412; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117222.4]
  assign _T_413 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117223.4]
  assign _T_414 = _T_413 | sectored_entries_6_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117224.4]
  assign _T_415 = _T_414 | sectored_entries_6_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117225.4]
  assign _T_416 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117226.4]
  assign _T_417 = _T_416[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117227.4]
  assign _T_418 = _T_417 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117228.4]
  assign sector_hits_6 = _T_415 & _T_418; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117229.4]
  assign _T_419 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117230.4]
  assign _T_420 = _T_419 | sectored_entries_7_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117231.4]
  assign _T_421 = _T_420 | sectored_entries_7_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@117232.4]
  assign _T_422 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@117233.4]
  assign _T_423 = _T_422[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@117234.4]
  assign _T_424 = _T_423 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@117235.4]
  assign sector_hits_7 = _T_421 & _T_424; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@117236.4]
  assign _T_427 = superpage_entries_0_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117239.4]
  assign _T_428 = vpn[19:10]; // @[TLB.scala 108:86:freechips.rocketchip.system.DefaultRV32Config.fir@117240.4]
  assign _T_429 = _T_427 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117241.4]
  assign superpage_hits_0 = superpage_entries_0_valid_0 & _T_429; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117243.4]
  assign _T_435 = vpn[9:0]; // @[TLB.scala 108:86:freechips.rocketchip.system.DefaultRV32Config.fir@117247.4]
  assign _T_440 = superpage_entries_1_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117253.4]
  assign _T_442 = _T_440 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117255.4]
  assign superpage_hits_1 = superpage_entries_1_valid_0 & _T_442; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117257.4]
  assign _T_453 = superpage_entries_2_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117267.4]
  assign _T_455 = _T_453 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117269.4]
  assign superpage_hits_2 = superpage_entries_2_valid_0 & _T_455; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117271.4]
  assign _T_466 = superpage_entries_3_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117281.4]
  assign _T_468 = _T_466 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117283.4]
  assign superpage_hits_3 = superpage_entries_3_valid_0 & _T_468; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117285.4]
  assign _T_477 = vpn[1:0]; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@117293.4]
  assign _GEN_1 = 2'h1 == _T_477 ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117297.4]
  assign _GEN_2 = 2'h2 == _T_477 ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117297.4]
  assign _GEN_3 = 2'h3 == _T_477 ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117297.4]
  assign _T_481 = _GEN_3 & _T_382; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117297.4]
  assign hitsVec_0 = vm_enabled & _T_481; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117298.4]
  assign _GEN_5 = 2'h1 == _T_477 ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117303.4]
  assign _GEN_6 = 2'h2 == _T_477 ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117303.4]
  assign _GEN_7 = 2'h3 == _T_477 ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117303.4]
  assign _T_486 = _GEN_7 & _T_388; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117303.4]
  assign hitsVec_1 = vm_enabled & _T_486; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117304.4]
  assign _GEN_9 = 2'h1 == _T_477 ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117309.4]
  assign _GEN_10 = 2'h2 == _T_477 ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117309.4]
  assign _GEN_11 = 2'h3 == _T_477 ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117309.4]
  assign _T_491 = _GEN_11 & _T_394; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117309.4]
  assign hitsVec_2 = vm_enabled & _T_491; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117310.4]
  assign _GEN_13 = 2'h1 == _T_477 ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117315.4]
  assign _GEN_14 = 2'h2 == _T_477 ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117315.4]
  assign _GEN_15 = 2'h3 == _T_477 ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117315.4]
  assign _T_496 = _GEN_15 & _T_400; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117315.4]
  assign hitsVec_3 = vm_enabled & _T_496; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117316.4]
  assign _GEN_17 = 2'h1 == _T_477 ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117321.4]
  assign _GEN_18 = 2'h2 == _T_477 ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117321.4]
  assign _GEN_19 = 2'h3 == _T_477 ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117321.4]
  assign _T_501 = _GEN_19 & _T_406; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117321.4]
  assign hitsVec_4 = vm_enabled & _T_501; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117322.4]
  assign _GEN_21 = 2'h1 == _T_477 ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117327.4]
  assign _GEN_22 = 2'h2 == _T_477 ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117327.4]
  assign _GEN_23 = 2'h3 == _T_477 ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117327.4]
  assign _T_506 = _GEN_23 & _T_412; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117327.4]
  assign hitsVec_5 = vm_enabled & _T_506; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117328.4]
  assign _GEN_25 = 2'h1 == _T_477 ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117333.4]
  assign _GEN_26 = 2'h2 == _T_477 ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117333.4]
  assign _GEN_27 = 2'h3 == _T_477 ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117333.4]
  assign _T_511 = _GEN_27 & _T_418; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117333.4]
  assign hitsVec_6 = vm_enabled & _T_511; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117334.4]
  assign _GEN_29 = 2'h1 == _T_477 ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117339.4]
  assign _GEN_30 = 2'h2 == _T_477 ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117339.4]
  assign _GEN_31 = 2'h3 == _T_477 ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117339.4]
  assign _T_516 = _GEN_31 & _T_424; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@117339.4]
  assign hitsVec_7 = vm_enabled & _T_516; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117340.4]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117355.4]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117370.4]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117385.4]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117400.4]
  assign _T_575 = special_entry_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117403.4]
  assign _T_577 = _T_575 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117405.4]
  assign _T_579 = special_entry_valid_0 & _T_577; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117407.4]
  assign _T_582 = special_entry_tag[9:0]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@117410.4]
  assign _T_584 = _T_582 == _T_435; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@117412.4]
  assign _T_585 = _T_25 | _T_584; // @[TLB.scala 108:42:freechips.rocketchip.system.DefaultRV32Config.fir@117413.4]
  assign _T_586 = _T_579 & _T_585; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@117414.4]
  assign hitsVec_12 = vm_enabled & _T_586; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@117415.4]
  assign _T_591 = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117420.4]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_591}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117427.4]
  assign _T_598 = vm_enabled == 1'h0; // @[TLB.scala 211:18:freechips.rocketchip.system.DefaultRV32Config.fir@117428.4]
  assign hits = {_T_598,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_591}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117429.4]
  assign _GEN_33 = 2'h1 == _T_477 ? sectored_entries_0_data_1 : sectored_entries_0_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117436.4]
  assign _GEN_34 = 2'h2 == _T_477 ? sectored_entries_0_data_2 : _GEN_33; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117436.4]
  assign _GEN_35 = 2'h3 == _T_477 ? sectored_entries_0_data_3 : _GEN_34; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117436.4]
  assign _GEN_37 = 2'h1 == _T_477 ? sectored_entries_1_data_1 : sectored_entries_1_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117477.4]
  assign _GEN_38 = 2'h2 == _T_477 ? sectored_entries_1_data_2 : _GEN_37; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117477.4]
  assign _GEN_39 = 2'h3 == _T_477 ? sectored_entries_1_data_3 : _GEN_38; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117477.4]
  assign _GEN_41 = 2'h1 == _T_477 ? sectored_entries_2_data_1 : sectored_entries_2_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117518.4]
  assign _GEN_42 = 2'h2 == _T_477 ? sectored_entries_2_data_2 : _GEN_41; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117518.4]
  assign _GEN_43 = 2'h3 == _T_477 ? sectored_entries_2_data_3 : _GEN_42; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117518.4]
  assign _GEN_45 = 2'h1 == _T_477 ? sectored_entries_3_data_1 : sectored_entries_3_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117559.4]
  assign _GEN_46 = 2'h2 == _T_477 ? sectored_entries_3_data_2 : _GEN_45; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117559.4]
  assign _GEN_47 = 2'h3 == _T_477 ? sectored_entries_3_data_3 : _GEN_46; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117559.4]
  assign _GEN_49 = 2'h1 == _T_477 ? sectored_entries_4_data_1 : sectored_entries_4_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117600.4]
  assign _GEN_50 = 2'h2 == _T_477 ? sectored_entries_4_data_2 : _GEN_49; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117600.4]
  assign _GEN_51 = 2'h3 == _T_477 ? sectored_entries_4_data_3 : _GEN_50; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117600.4]
  assign _GEN_53 = 2'h1 == _T_477 ? sectored_entries_5_data_1 : sectored_entries_5_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117641.4]
  assign _GEN_54 = 2'h2 == _T_477 ? sectored_entries_5_data_2 : _GEN_53; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117641.4]
  assign _GEN_55 = 2'h3 == _T_477 ? sectored_entries_5_data_3 : _GEN_54; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117641.4]
  assign _GEN_57 = 2'h1 == _T_477 ? sectored_entries_6_data_1 : sectored_entries_6_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117682.4]
  assign _GEN_58 = 2'h2 == _T_477 ? sectored_entries_6_data_2 : _GEN_57; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117682.4]
  assign _GEN_59 = 2'h3 == _T_477 ? sectored_entries_6_data_3 : _GEN_58; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117682.4]
  assign _GEN_61 = 2'h1 == _T_477 ? sectored_entries_7_data_1 : sectored_entries_7_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117723.4]
  assign _GEN_62 = 2'h2 == _T_477 ? sectored_entries_7_data_2 : _GEN_61; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117723.4]
  assign _GEN_63 = 2'h3 == _T_477 ? sectored_entries_7_data_3 : _GEN_62; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@117723.4]
  assign _T_758 = superpage_entries_0_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@117788.4]
  assign _T_761 = _2_9_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117799.4]
  assign _T_765 = vpn | _2_9_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117803.4]
  assign _T_766 = _T_765[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117804.4]
  assign _T_767 = {_T_761,_T_766}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117805.4]
  assign _T_782 = superpage_entries_1_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@117835.4]
  assign _T_785 = _2_10_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117846.4]
  assign _T_789 = vpn | _2_10_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117850.4]
  assign _T_790 = _T_789[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117851.4]
  assign _T_791 = {_T_785,_T_790}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117852.4]
  assign _T_806 = superpage_entries_2_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@117882.4]
  assign _T_809 = _2_11_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117893.4]
  assign _T_813 = vpn | _2_11_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117897.4]
  assign _T_814 = _T_813[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117898.4]
  assign _T_815 = {_T_809,_T_814}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117899.4]
  assign _T_830 = superpage_entries_3_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@117929.4]
  assign _T_833 = _2_12_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117940.4]
  assign _T_837 = vpn | _2_12_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117944.4]
  assign _T_838 = _T_837[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117945.4]
  assign _T_839 = {_T_833,_T_838}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117946.4]
  assign _T_857 = _2_13_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@117987.4]
  assign _T_861 = _T_27 | _2_13_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@117991.4]
  assign _T_862 = _T_861[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@117992.4]
  assign _T_863 = {_T_857,_T_862}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@117993.4]
  assign _T_865 = hitsVec_0 ? _2_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117995.4]
  assign _T_866 = hitsVec_1 ? _2_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117996.4]
  assign _T_867 = hitsVec_2 ? _2_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117997.4]
  assign _T_868 = hitsVec_3 ? _2_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117998.4]
  assign _T_869 = hitsVec_4 ? _2_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@117999.4]
  assign _T_870 = hitsVec_5 ? _2_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118000.4]
  assign _T_871 = hitsVec_6 ? _2_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118001.4]
  assign _T_872 = hitsVec_7 ? _2_8_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118002.4]
  assign _T_873 = hitsVec_8 ? _T_767 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118003.4]
  assign _T_874 = hitsVec_9 ? _T_791 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118004.4]
  assign _T_875 = hitsVec_10 ? _T_815 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118005.4]
  assign _T_876 = hitsVec_11 ? _T_839 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118006.4]
  assign _T_877 = hitsVec_12 ? _T_863 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118007.4]
  assign _T_878 = _T_598 ? vpn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118008.4]
  assign _T_879 = _T_865 | _T_866; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118009.4]
  assign _T_880 = _T_879 | _T_867; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118010.4]
  assign _T_881 = _T_880 | _T_868; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118011.4]
  assign _T_882 = _T_881 | _T_869; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118012.4]
  assign _T_883 = _T_882 | _T_870; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118013.4]
  assign _T_884 = _T_883 | _T_871; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118014.4]
  assign _T_885 = _T_884 | _T_872; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118015.4]
  assign _T_886 = _T_885 | _T_873; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118016.4]
  assign _T_887 = _T_886 | _T_874; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118017.4]
  assign _T_888 = _T_887 | _T_875; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118018.4]
  assign _T_889 = _T_888 | _T_876; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118019.4]
  assign _T_890 = _T_889 | _T_877; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118020.4]
  assign ppn = _T_890 | _T_878; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@118021.4]
  assign _T_892 = invalidate_refill == 1'h0; // @[TLB.scala 215:22:freechips.rocketchip.system.DefaultRV32Config.fir@118024.4]
  assign _T_893 = io_ptw_resp_valid & _T_892; // @[TLB.scala 215:19:freechips.rocketchip.system.DefaultRV32Config.fir@118025.4]
  assign _T_895 = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 221:25:freechips.rocketchip.system.DefaultRV32Config.fir@118032.6]
  assign _T_896 = io_ptw_resp_bits_pte_w == 1'h0; // @[PTW.scala 68:47:freechips.rocketchip.system.DefaultRV32Config.fir@118035.6]
  assign _T_897 = io_ptw_resp_bits_pte_x & _T_896; // @[PTW.scala 68:44:freechips.rocketchip.system.DefaultRV32Config.fir@118036.6]
  assign _T_898 = io_ptw_resp_bits_pte_r | _T_897; // @[PTW.scala 68:38:freechips.rocketchip.system.DefaultRV32Config.fir@118037.6]
  assign _T_899 = io_ptw_resp_bits_pte_v & _T_898; // @[PTW.scala 68:32:freechips.rocketchip.system.DefaultRV32Config.fir@118038.6]
  assign _T_900 = _T_899 & io_ptw_resp_bits_pte_a; // @[PTW.scala 68:52:freechips.rocketchip.system.DefaultRV32Config.fir@118039.6]
  assign _T_901 = _T_900 & io_ptw_resp_bits_pte_r; // @[PTW.scala 72:35:freechips.rocketchip.system.DefaultRV32Config.fir@118040.6]
  assign _T_907 = _T_900 & io_ptw_resp_bits_pte_w; // @[PTW.scala 73:35:freechips.rocketchip.system.DefaultRV32Config.fir@118047.6]
  assign _T_908 = _T_907 & io_ptw_resp_bits_pte_d; // @[PTW.scala 73:40:freechips.rocketchip.system.DefaultRV32Config.fir@118048.6]
  assign _T_914 = _T_900 & io_ptw_resp_bits_pte_x; // @[PTW.scala 74:35:freechips.rocketchip.system.DefaultRV32Config.fir@118055.6]
  assign _T_915 = io_ptw_resp_bits_homogeneous == 1'h0; // @[TLB.scala 234:37:freechips.rocketchip.system.DefaultRV32Config.fir@118064.6]
  assign _T_923 = {prot_x,prot_r,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 136:26:freechips.rocketchip.system.DefaultRV32Config.fir@118076.8]
  assign _T_931 = {refill_ppn,io_ptw_resp_bits_pte_u,_T_895,io_ptw_resp_bits_ae,_T_908,_T_914,_T_901,prot_w,_T_923}; // @[TLB.scala 136:26:freechips.rocketchip.system.DefaultRV32Config.fir@118084.8]
  assign _T_932 = io_ptw_resp_bits_level < 1'h1; // @[TLB.scala 236:40:freechips.rocketchip.system.DefaultRV32Config.fir@118088.8]
  assign _T_933 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@118090.10]
  assign _GEN_66 = _T_933 | superpage_entries_0_valid_0; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@118091.10]
  assign _T_948 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@118111.10]
  assign _GEN_70 = _T_948 | superpage_entries_1_valid_0; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@118112.10]
  assign _T_963 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@118132.10]
  assign _GEN_74 = _T_963 | superpage_entries_2_valid_0; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@118133.10]
  assign _T_978 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@118153.10]
  assign _GEN_78 = _T_978 | superpage_entries_3_valid_0; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@118154.10]
  assign _T_993 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 241:22:freechips.rocketchip.system.DefaultRV32Config.fir@118176.10]
  assign _T_994 = _T_993 == 3'h0; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118177.10]
  assign _T_995 = r_sectored_hit == 1'h0; // @[TLB.scala 243:15:freechips.rocketchip.system.DefaultRV32Config.fir@118179.12]
  assign _GEN_80 = _T_995 ? 1'h0 : sectored_entries_0_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118180.12]
  assign _GEN_81 = _T_995 ? 1'h0 : sectored_entries_0_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118180.12]
  assign _GEN_82 = _T_995 ? 1'h0 : sectored_entries_0_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118180.12]
  assign _GEN_83 = _T_995 ? 1'h0 : sectored_entries_0_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118180.12]
  assign _T_996 = r_refill_tag[1:0]; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@118188.12]
  assign _GEN_950 = 2'h0 == _T_996; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  assign _GEN_84 = _GEN_950 | _GEN_80; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  assign _GEN_951 = 2'h1 == _T_996; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  assign _GEN_85 = _GEN_951 | _GEN_81; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  assign _GEN_952 = 2'h2 == _T_996; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  assign _GEN_86 = _GEN_952 | _GEN_82; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  assign _GEN_953 = 2'h3 == _T_996; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  assign _GEN_87 = _GEN_953 | _GEN_83; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118189.12]
  assign _GEN_92 = _T_994 ? _GEN_84 : sectored_entries_0_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118178.10]
  assign _GEN_93 = _T_994 ? _GEN_85 : sectored_entries_0_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118178.10]
  assign _GEN_94 = _T_994 ? _GEN_86 : sectored_entries_0_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118178.10]
  assign _GEN_95 = _T_994 ? _GEN_87 : sectored_entries_0_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118178.10]
  assign _T_1011 = _T_993 == 3'h1; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118206.10]
  assign _GEN_102 = _T_995 ? 1'h0 : sectored_entries_1_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118209.12]
  assign _GEN_103 = _T_995 ? 1'h0 : sectored_entries_1_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118209.12]
  assign _GEN_104 = _T_995 ? 1'h0 : sectored_entries_1_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118209.12]
  assign _GEN_105 = _T_995 ? 1'h0 : sectored_entries_1_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118209.12]
  assign _GEN_106 = _GEN_950 | _GEN_102; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118218.12]
  assign _GEN_107 = _GEN_951 | _GEN_103; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118218.12]
  assign _GEN_108 = _GEN_952 | _GEN_104; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118218.12]
  assign _GEN_109 = _GEN_953 | _GEN_105; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118218.12]
  assign _GEN_114 = _T_1011 ? _GEN_106 : sectored_entries_1_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118207.10]
  assign _GEN_115 = _T_1011 ? _GEN_107 : sectored_entries_1_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118207.10]
  assign _GEN_116 = _T_1011 ? _GEN_108 : sectored_entries_1_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118207.10]
  assign _GEN_117 = _T_1011 ? _GEN_109 : sectored_entries_1_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118207.10]
  assign _T_1028 = _T_993 == 3'h2; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118235.10]
  assign _GEN_124 = _T_995 ? 1'h0 : sectored_entries_2_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118238.12]
  assign _GEN_125 = _T_995 ? 1'h0 : sectored_entries_2_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118238.12]
  assign _GEN_126 = _T_995 ? 1'h0 : sectored_entries_2_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118238.12]
  assign _GEN_127 = _T_995 ? 1'h0 : sectored_entries_2_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118238.12]
  assign _GEN_128 = _GEN_950 | _GEN_124; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118247.12]
  assign _GEN_129 = _GEN_951 | _GEN_125; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118247.12]
  assign _GEN_130 = _GEN_952 | _GEN_126; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118247.12]
  assign _GEN_131 = _GEN_953 | _GEN_127; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118247.12]
  assign _GEN_136 = _T_1028 ? _GEN_128 : sectored_entries_2_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118236.10]
  assign _GEN_137 = _T_1028 ? _GEN_129 : sectored_entries_2_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118236.10]
  assign _GEN_138 = _T_1028 ? _GEN_130 : sectored_entries_2_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118236.10]
  assign _GEN_139 = _T_1028 ? _GEN_131 : sectored_entries_2_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118236.10]
  assign _T_1045 = _T_993 == 3'h3; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118264.10]
  assign _GEN_146 = _T_995 ? 1'h0 : sectored_entries_3_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118267.12]
  assign _GEN_147 = _T_995 ? 1'h0 : sectored_entries_3_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118267.12]
  assign _GEN_148 = _T_995 ? 1'h0 : sectored_entries_3_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118267.12]
  assign _GEN_149 = _T_995 ? 1'h0 : sectored_entries_3_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118267.12]
  assign _GEN_150 = _GEN_950 | _GEN_146; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118276.12]
  assign _GEN_151 = _GEN_951 | _GEN_147; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118276.12]
  assign _GEN_152 = _GEN_952 | _GEN_148; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118276.12]
  assign _GEN_153 = _GEN_953 | _GEN_149; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118276.12]
  assign _GEN_158 = _T_1045 ? _GEN_150 : sectored_entries_3_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118265.10]
  assign _GEN_159 = _T_1045 ? _GEN_151 : sectored_entries_3_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118265.10]
  assign _GEN_160 = _T_1045 ? _GEN_152 : sectored_entries_3_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118265.10]
  assign _GEN_161 = _T_1045 ? _GEN_153 : sectored_entries_3_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118265.10]
  assign _T_1062 = _T_993 == 3'h4; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118293.10]
  assign _GEN_168 = _T_995 ? 1'h0 : sectored_entries_4_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118296.12]
  assign _GEN_169 = _T_995 ? 1'h0 : sectored_entries_4_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118296.12]
  assign _GEN_170 = _T_995 ? 1'h0 : sectored_entries_4_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118296.12]
  assign _GEN_171 = _T_995 ? 1'h0 : sectored_entries_4_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118296.12]
  assign _GEN_172 = _GEN_950 | _GEN_168; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118305.12]
  assign _GEN_173 = _GEN_951 | _GEN_169; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118305.12]
  assign _GEN_174 = _GEN_952 | _GEN_170; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118305.12]
  assign _GEN_175 = _GEN_953 | _GEN_171; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118305.12]
  assign _GEN_180 = _T_1062 ? _GEN_172 : sectored_entries_4_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118294.10]
  assign _GEN_181 = _T_1062 ? _GEN_173 : sectored_entries_4_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118294.10]
  assign _GEN_182 = _T_1062 ? _GEN_174 : sectored_entries_4_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118294.10]
  assign _GEN_183 = _T_1062 ? _GEN_175 : sectored_entries_4_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118294.10]
  assign _T_1079 = _T_993 == 3'h5; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118322.10]
  assign _GEN_190 = _T_995 ? 1'h0 : sectored_entries_5_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118325.12]
  assign _GEN_191 = _T_995 ? 1'h0 : sectored_entries_5_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118325.12]
  assign _GEN_192 = _T_995 ? 1'h0 : sectored_entries_5_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118325.12]
  assign _GEN_193 = _T_995 ? 1'h0 : sectored_entries_5_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118325.12]
  assign _GEN_194 = _GEN_950 | _GEN_190; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118334.12]
  assign _GEN_195 = _GEN_951 | _GEN_191; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118334.12]
  assign _GEN_196 = _GEN_952 | _GEN_192; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118334.12]
  assign _GEN_197 = _GEN_953 | _GEN_193; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118334.12]
  assign _GEN_202 = _T_1079 ? _GEN_194 : sectored_entries_5_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118323.10]
  assign _GEN_203 = _T_1079 ? _GEN_195 : sectored_entries_5_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118323.10]
  assign _GEN_204 = _T_1079 ? _GEN_196 : sectored_entries_5_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118323.10]
  assign _GEN_205 = _T_1079 ? _GEN_197 : sectored_entries_5_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118323.10]
  assign _T_1096 = _T_993 == 3'h6; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118351.10]
  assign _GEN_212 = _T_995 ? 1'h0 : sectored_entries_6_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118354.12]
  assign _GEN_213 = _T_995 ? 1'h0 : sectored_entries_6_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118354.12]
  assign _GEN_214 = _T_995 ? 1'h0 : sectored_entries_6_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118354.12]
  assign _GEN_215 = _T_995 ? 1'h0 : sectored_entries_6_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118354.12]
  assign _GEN_216 = _GEN_950 | _GEN_212; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118363.12]
  assign _GEN_217 = _GEN_951 | _GEN_213; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118363.12]
  assign _GEN_218 = _GEN_952 | _GEN_214; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118363.12]
  assign _GEN_219 = _GEN_953 | _GEN_215; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118363.12]
  assign _GEN_224 = _T_1096 ? _GEN_216 : sectored_entries_6_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118352.10]
  assign _GEN_225 = _T_1096 ? _GEN_217 : sectored_entries_6_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118352.10]
  assign _GEN_226 = _T_1096 ? _GEN_218 : sectored_entries_6_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118352.10]
  assign _GEN_227 = _T_1096 ? _GEN_219 : sectored_entries_6_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118352.10]
  assign _T_1113 = _T_993 == 3'h7; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@118380.10]
  assign _GEN_234 = _T_995 ? 1'h0 : sectored_entries_7_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118383.12]
  assign _GEN_235 = _T_995 ? 1'h0 : sectored_entries_7_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118383.12]
  assign _GEN_236 = _T_995 ? 1'h0 : sectored_entries_7_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118383.12]
  assign _GEN_237 = _T_995 ? 1'h0 : sectored_entries_7_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@118383.12]
  assign _GEN_238 = _GEN_950 | _GEN_234; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118392.12]
  assign _GEN_239 = _GEN_951 | _GEN_235; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118392.12]
  assign _GEN_240 = _GEN_952 | _GEN_236; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118392.12]
  assign _GEN_241 = _GEN_953 | _GEN_237; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@118392.12]
  assign _GEN_246 = _T_1113 ? _GEN_238 : sectored_entries_7_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118381.10]
  assign _GEN_247 = _T_1113 ? _GEN_239 : sectored_entries_7_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118381.10]
  assign _GEN_248 = _T_1113 ? _GEN_240 : sectored_entries_7_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118381.10]
  assign _GEN_249 = _T_1113 ? _GEN_241 : sectored_entries_7_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@118381.10]
  assign _GEN_258 = _T_932 ? _GEN_66 : superpage_entries_0_valid_0; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_262 = _T_932 ? _GEN_70 : superpage_entries_1_valid_0; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_266 = _T_932 ? _GEN_74 : superpage_entries_2_valid_0; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_270 = _T_932 ? _GEN_78 : superpage_entries_3_valid_0; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_272 = _T_932 ? sectored_entries_0_valid_0 : _GEN_92; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_273 = _T_932 ? sectored_entries_0_valid_1 : _GEN_93; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_274 = _T_932 ? sectored_entries_0_valid_2 : _GEN_94; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_275 = _T_932 ? sectored_entries_0_valid_3 : _GEN_95; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_282 = _T_932 ? sectored_entries_1_valid_0 : _GEN_114; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_283 = _T_932 ? sectored_entries_1_valid_1 : _GEN_115; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_284 = _T_932 ? sectored_entries_1_valid_2 : _GEN_116; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_285 = _T_932 ? sectored_entries_1_valid_3 : _GEN_117; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_292 = _T_932 ? sectored_entries_2_valid_0 : _GEN_136; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_293 = _T_932 ? sectored_entries_2_valid_1 : _GEN_137; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_294 = _T_932 ? sectored_entries_2_valid_2 : _GEN_138; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_295 = _T_932 ? sectored_entries_2_valid_3 : _GEN_139; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_302 = _T_932 ? sectored_entries_3_valid_0 : _GEN_158; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_303 = _T_932 ? sectored_entries_3_valid_1 : _GEN_159; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_304 = _T_932 ? sectored_entries_3_valid_2 : _GEN_160; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_305 = _T_932 ? sectored_entries_3_valid_3 : _GEN_161; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_312 = _T_932 ? sectored_entries_4_valid_0 : _GEN_180; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_313 = _T_932 ? sectored_entries_4_valid_1 : _GEN_181; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_314 = _T_932 ? sectored_entries_4_valid_2 : _GEN_182; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_315 = _T_932 ? sectored_entries_4_valid_3 : _GEN_183; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_322 = _T_932 ? sectored_entries_5_valid_0 : _GEN_202; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_323 = _T_932 ? sectored_entries_5_valid_1 : _GEN_203; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_324 = _T_932 ? sectored_entries_5_valid_2 : _GEN_204; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_325 = _T_932 ? sectored_entries_5_valid_3 : _GEN_205; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_332 = _T_932 ? sectored_entries_6_valid_0 : _GEN_224; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_333 = _T_932 ? sectored_entries_6_valid_1 : _GEN_225; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_334 = _T_932 ? sectored_entries_6_valid_2 : _GEN_226; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_335 = _T_932 ? sectored_entries_6_valid_3 : _GEN_227; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_342 = _T_932 ? sectored_entries_7_valid_0 : _GEN_246; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_343 = _T_932 ? sectored_entries_7_valid_1 : _GEN_247; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_344 = _T_932 ? sectored_entries_7_valid_2 : _GEN_248; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_345 = _T_932 ? sectored_entries_7_valid_3 : _GEN_249; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@118089.8]
  assign _GEN_354 = _T_915 | special_entry_valid_0; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_358 = _T_915 ? superpage_entries_0_valid_0 : _GEN_258; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_362 = _T_915 ? superpage_entries_1_valid_0 : _GEN_262; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_366 = _T_915 ? superpage_entries_2_valid_0 : _GEN_266; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_370 = _T_915 ? superpage_entries_3_valid_0 : _GEN_270; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_372 = _T_915 ? sectored_entries_0_valid_0 : _GEN_272; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_373 = _T_915 ? sectored_entries_0_valid_1 : _GEN_273; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_374 = _T_915 ? sectored_entries_0_valid_2 : _GEN_274; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_375 = _T_915 ? sectored_entries_0_valid_3 : _GEN_275; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_382 = _T_915 ? sectored_entries_1_valid_0 : _GEN_282; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_383 = _T_915 ? sectored_entries_1_valid_1 : _GEN_283; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_384 = _T_915 ? sectored_entries_1_valid_2 : _GEN_284; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_385 = _T_915 ? sectored_entries_1_valid_3 : _GEN_285; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_392 = _T_915 ? sectored_entries_2_valid_0 : _GEN_292; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_393 = _T_915 ? sectored_entries_2_valid_1 : _GEN_293; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_394 = _T_915 ? sectored_entries_2_valid_2 : _GEN_294; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_395 = _T_915 ? sectored_entries_2_valid_3 : _GEN_295; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_402 = _T_915 ? sectored_entries_3_valid_0 : _GEN_302; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_403 = _T_915 ? sectored_entries_3_valid_1 : _GEN_303; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_404 = _T_915 ? sectored_entries_3_valid_2 : _GEN_304; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_405 = _T_915 ? sectored_entries_3_valid_3 : _GEN_305; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_412 = _T_915 ? sectored_entries_4_valid_0 : _GEN_312; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_413 = _T_915 ? sectored_entries_4_valid_1 : _GEN_313; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_414 = _T_915 ? sectored_entries_4_valid_2 : _GEN_314; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_415 = _T_915 ? sectored_entries_4_valid_3 : _GEN_315; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_422 = _T_915 ? sectored_entries_5_valid_0 : _GEN_322; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_423 = _T_915 ? sectored_entries_5_valid_1 : _GEN_323; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_424 = _T_915 ? sectored_entries_5_valid_2 : _GEN_324; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_425 = _T_915 ? sectored_entries_5_valid_3 : _GEN_325; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_432 = _T_915 ? sectored_entries_6_valid_0 : _GEN_332; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_433 = _T_915 ? sectored_entries_6_valid_1 : _GEN_333; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_434 = _T_915 ? sectored_entries_6_valid_2 : _GEN_334; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_435 = _T_915 ? sectored_entries_6_valid_3 : _GEN_335; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_442 = _T_915 ? sectored_entries_7_valid_0 : _GEN_342; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_443 = _T_915 ? sectored_entries_7_valid_1 : _GEN_343; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_444 = _T_915 ? sectored_entries_7_valid_2 : _GEN_344; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_445 = _T_915 ? sectored_entries_7_valid_3 : _GEN_345; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@118066.6]
  assign _GEN_454 = _T_893 ? _GEN_354 : special_entry_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_458 = _T_893 ? _GEN_358 : superpage_entries_0_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_462 = _T_893 ? _GEN_362 : superpage_entries_1_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_466 = _T_893 ? _GEN_366 : superpage_entries_2_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_470 = _T_893 ? _GEN_370 : superpage_entries_3_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_472 = _T_893 ? _GEN_372 : sectored_entries_0_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_473 = _T_893 ? _GEN_373 : sectored_entries_0_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_474 = _T_893 ? _GEN_374 : sectored_entries_0_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_475 = _T_893 ? _GEN_375 : sectored_entries_0_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_482 = _T_893 ? _GEN_382 : sectored_entries_1_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_483 = _T_893 ? _GEN_383 : sectored_entries_1_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_484 = _T_893 ? _GEN_384 : sectored_entries_1_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_485 = _T_893 ? _GEN_385 : sectored_entries_1_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_492 = _T_893 ? _GEN_392 : sectored_entries_2_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_493 = _T_893 ? _GEN_393 : sectored_entries_2_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_494 = _T_893 ? _GEN_394 : sectored_entries_2_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_495 = _T_893 ? _GEN_395 : sectored_entries_2_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_502 = _T_893 ? _GEN_402 : sectored_entries_3_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_503 = _T_893 ? _GEN_403 : sectored_entries_3_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_504 = _T_893 ? _GEN_404 : sectored_entries_3_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_505 = _T_893 ? _GEN_405 : sectored_entries_3_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_512 = _T_893 ? _GEN_412 : sectored_entries_4_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_513 = _T_893 ? _GEN_413 : sectored_entries_4_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_514 = _T_893 ? _GEN_414 : sectored_entries_4_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_515 = _T_893 ? _GEN_415 : sectored_entries_4_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_522 = _T_893 ? _GEN_422 : sectored_entries_5_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_523 = _T_893 ? _GEN_423 : sectored_entries_5_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_524 = _T_893 ? _GEN_424 : sectored_entries_5_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_525 = _T_893 ? _GEN_425 : sectored_entries_5_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_532 = _T_893 ? _GEN_432 : sectored_entries_6_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_533 = _T_893 ? _GEN_433 : sectored_entries_6_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_534 = _T_893 ? _GEN_434 : sectored_entries_6_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_535 = _T_893 ? _GEN_435 : sectored_entries_6_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_542 = _T_893 ? _GEN_442 : sectored_entries_7_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_543 = _T_893 ? _GEN_443 : sectored_entries_7_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_544 = _T_893 ? _GEN_444 : sectored_entries_7_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _GEN_545 = _T_893 ? _GEN_445 : sectored_entries_7_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@118026.4]
  assign _T_1575 = {_2_19_io_y_ae,_2_18_io_y_ae,_2_17_io_y_ae,_2_16_io_y_ae,_2_15_io_y_ae,_2_14_io_y_ae}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119431.4]
  assign ptw_ae_array = {1'h0,_2_26_io_y_ae,_2_25_io_y_ae,_2_24_io_y_ae,_2_23_io_y_ae,_2_22_io_y_ae,_2_21_io_y_ae,_2_20_io_y_ae,_T_1575}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119439.4]
  assign _T_1583 = priv_s == 1'h0; // @[TLB.scala 253:24:freechips.rocketchip.system.DefaultRV32Config.fir@119440.4]
  assign _T_1584 = _T_1583 | io_ptw_status_sum; // @[TLB.scala 253:32:freechips.rocketchip.system.DefaultRV32Config.fir@119441.4]
  assign _T_1589 = {_2_19_io_y_u,_2_18_io_y_u,_2_17_io_y_u,_2_16_io_y_u,_2_15_io_y_u,_2_14_io_y_u}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119446.4]
  assign _T_1596 = {_2_26_io_y_u,_2_25_io_y_u,_2_24_io_y_u,_2_23_io_y_u,_2_22_io_y_u,_2_21_io_y_u,_2_20_io_y_u,_T_1589}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119453.4]
  assign _T_1597 = _T_1584 ? _T_1596 : 13'h0; // @[TLB.scala 253:23:freechips.rocketchip.system.DefaultRV32Config.fir@119454.4]
  assign _T_1610 = ~ _T_1596; // @[TLB.scala 253:98:freechips.rocketchip.system.DefaultRV32Config.fir@119467.4]
  assign _T_1611 = priv_s ? _T_1610 : 13'h0; // @[TLB.scala 253:89:freechips.rocketchip.system.DefaultRV32Config.fir@119468.4]
  assign priv_rw_ok = _T_1597 | _T_1611; // @[TLB.scala 253:84:freechips.rocketchip.system.DefaultRV32Config.fir@119469.4]
  assign _T_1641 = {_2_19_io_y_sr,_2_18_io_y_sr,_2_17_io_y_sr,_2_16_io_y_sr,_2_15_io_y_sr,_2_14_io_y_sr}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119500.4]
  assign _T_1648 = {_2_26_io_y_sr,_2_25_io_y_sr,_2_24_io_y_sr,_2_23_io_y_sr,_2_22_io_y_sr,_2_21_io_y_sr,_2_20_io_y_sr,_T_1641}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119507.4]
  assign _T_1653 = {_2_19_io_y_sx,_2_18_io_y_sx,_2_17_io_y_sx,_2_16_io_y_sx,_2_15_io_y_sx,_2_14_io_y_sx}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119512.4]
  assign _T_1660 = {_2_26_io_y_sx,_2_25_io_y_sx,_2_24_io_y_sx,_2_23_io_y_sx,_2_22_io_y_sx,_2_21_io_y_sx,_2_20_io_y_sx,_T_1653}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119519.4]
  assign _T_1661 = io_ptw_status_mxr ? _T_1660 : 13'h0; // @[TLB.scala 255:73:freechips.rocketchip.system.DefaultRV32Config.fir@119520.4]
  assign _T_1662 = _T_1648 | _T_1661; // @[TLB.scala 255:68:freechips.rocketchip.system.DefaultRV32Config.fir@119521.4]
  assign _T_1663 = priv_rw_ok & _T_1662; // @[TLB.scala 255:40:freechips.rocketchip.system.DefaultRV32Config.fir@119522.4]
  assign r_array = {1'h1,_T_1663}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119523.4]
  assign _T_1668 = {_2_19_io_y_sw,_2_18_io_y_sw,_2_17_io_y_sw,_2_16_io_y_sw,_2_15_io_y_sw,_2_14_io_y_sw}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119528.4]
  assign _T_1675 = {_2_26_io_y_sw,_2_25_io_y_sw,_2_24_io_y_sw,_2_23_io_y_sw,_2_22_io_y_sw,_2_21_io_y_sw,_2_20_io_y_sw,_T_1668}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119535.4]
  assign _T_1676 = priv_rw_ok & _T_1675; // @[TLB.scala 256:40:freechips.rocketchip.system.DefaultRV32Config.fir@119536.4]
  assign w_array = {1'h1,_T_1676}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119537.4]
  assign _T_1691 = prot_r ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119553.4]
  assign _T_1696 = {_2_32_io_y_pr,_2_31_io_y_pr,_2_30_io_y_pr,_2_29_io_y_pr,_2_28_io_y_pr,_2_27_io_y_pr}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119558.4]
  assign _T_1703 = {_T_1691,_2_38_io_y_pr,_2_37_io_y_pr,_2_36_io_y_pr,_2_35_io_y_pr,_2_34_io_y_pr,_2_33_io_y_pr,_T_1696}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119565.4]
  assign _T_1704 = ~ ptw_ae_array; // @[TLB.scala 258:89:freechips.rocketchip.system.DefaultRV32Config.fir@119566.4]
  assign pr_array = _T_1703 & _T_1704; // @[TLB.scala 258:87:freechips.rocketchip.system.DefaultRV32Config.fir@119567.4]
  assign _T_1706 = prot_w ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119569.4]
  assign _T_1711 = {_2_32_io_y_pw,_2_31_io_y_pw,_2_30_io_y_pw,_2_29_io_y_pw,_2_28_io_y_pw,_2_27_io_y_pw}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119574.4]
  assign _T_1718 = {_T_1706,_2_38_io_y_pw,_2_37_io_y_pw,_2_36_io_y_pw,_2_35_io_y_pw,_2_34_io_y_pw,_2_33_io_y_pw,_T_1711}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119581.4]
  assign pw_array = _T_1718 & _T_1704; // @[TLB.scala 259:87:freechips.rocketchip.system.DefaultRV32Config.fir@119583.4]
  assign _T_1736 = prot_eff ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119601.4]
  assign _T_1741 = {_2_32_io_y_eff,_2_31_io_y_eff,_2_30_io_y_eff,_2_29_io_y_eff,_2_28_io_y_eff,_2_27_io_y_eff}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119606.4]
  assign eff_array = {_T_1736,_2_38_io_y_eff,_2_37_io_y_eff,_2_36_io_y_eff,_2_35_io_y_eff,_2_34_io_y_eff,_2_33_io_y_eff,_T_1741}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119613.4]
  assign _T_1749 = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119615.4]
  assign _T_1754 = {_2_32_io_y_c,_2_31_io_y_c,_2_30_io_y_c,_2_29_io_y_c,_2_28_io_y_c,_2_27_io_y_c}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119620.4]
  assign c_array = {_T_1749,_2_38_io_y_c,_2_37_io_y_c,_2_36_io_y_c,_2_35_io_y_c,_2_34_io_y_c,_2_33_io_y_c,_T_1754}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119627.4]
  assign _T_1762 = prot_al ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@119629.4]
  assign _T_1767 = {_2_32_io_y_paa,_2_31_io_y_paa,_2_30_io_y_paa,_2_29_io_y_paa,_2_28_io_y_paa,_2_27_io_y_paa}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119634.4]
  assign paa_array = {_T_1762,_2_38_io_y_paa,_2_37_io_y_paa,_2_36_io_y_paa,_2_35_io_y_paa,_2_34_io_y_paa,_2_33_io_y_paa,_T_1767}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119641.4]
  assign _T_1780 = {_2_32_io_y_pal,_2_31_io_y_pal,_2_30_io_y_pal,_2_29_io_y_pal,_2_28_io_y_pal,_2_27_io_y_pal}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119648.4]
  assign pal_array = {_T_1762,_2_38_io_y_pal,_2_37_io_y_pal,_2_36_io_y_pal,_2_35_io_y_pal,_2_34_io_y_pal,_2_33_io_y_pal,_T_1780}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119655.4]
  assign paa_array_if_cached = paa_array | c_array; // @[TLB.scala 265:39:freechips.rocketchip.system.DefaultRV32Config.fir@119657.4]
  assign pal_array_if_cached = pal_array | c_array; // @[TLB.scala 266:39:freechips.rocketchip.system.DefaultRV32Config.fir@119659.4]
  assign _T_1802 = 4'h1 << io_req_bits_size; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@119674.4]
  assign _T_1804 = _T_1802 - 4'h1; // @[TLB.scala 269:69:freechips.rocketchip.system.DefaultRV32Config.fir@119676.4]
  assign _GEN_982 = {{28'd0}, _T_1804}; // @[TLB.scala 269:39:freechips.rocketchip.system.DefaultRV32Config.fir@119677.4]
  assign _T_1805 = io_req_bits_vaddr & _GEN_982; // @[TLB.scala 269:39:freechips.rocketchip.system.DefaultRV32Config.fir@119677.4]
  assign misaligned = _T_1805 != 32'h0; // @[TLB.scala 269:75:freechips.rocketchip.system.DefaultRV32Config.fir@119678.4]
  assign _T_1806 = io_req_bits_cmd == 5'h6; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119679.4]
  assign _T_1807 = io_req_bits_cmd == 5'h7; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119680.4]
  assign cmd_lrsc = _T_1806 | _T_1807; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119681.4]
  assign _T_1809 = io_req_bits_cmd == 5'h4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119683.4]
  assign _T_1810 = io_req_bits_cmd == 5'h9; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119684.4]
  assign _T_1811 = io_req_bits_cmd == 5'ha; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119685.4]
  assign _T_1812 = io_req_bits_cmd == 5'hb; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119686.4]
  assign _T_1813 = _T_1809 | _T_1810; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119687.4]
  assign _T_1814 = _T_1813 | _T_1811; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119688.4]
  assign cmd_amo_logical = _T_1814 | _T_1812; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119689.4]
  assign _T_1816 = io_req_bits_cmd == 5'h8; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119691.4]
  assign _T_1817 = io_req_bits_cmd == 5'hc; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119692.4]
  assign _T_1818 = io_req_bits_cmd == 5'hd; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119693.4]
  assign _T_1819 = io_req_bits_cmd == 5'he; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119694.4]
  assign _T_1820 = io_req_bits_cmd == 5'hf; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119695.4]
  assign _T_1821 = _T_1816 | _T_1817; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119696.4]
  assign _T_1822 = _T_1821 | _T_1818; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119697.4]
  assign _T_1823 = _T_1822 | _T_1819; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119698.4]
  assign cmd_amo_arithmetic = _T_1823 | _T_1820; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119699.4]
  assign _T_1825 = io_req_bits_cmd == 5'h0; // @[Consts.scala 82:31:freechips.rocketchip.system.DefaultRV32Config.fir@119701.4]
  assign _T_1827 = _T_1825 | _T_1806; // @[Consts.scala 82:41:freechips.rocketchip.system.DefaultRV32Config.fir@119703.4]
  assign _T_1829 = _T_1827 | _T_1807; // @[Consts.scala 82:58:freechips.rocketchip.system.DefaultRV32Config.fir@119705.4]
  assign _T_1846 = cmd_amo_logical | cmd_amo_arithmetic; // @[Consts.scala 80:44:freechips.rocketchip.system.DefaultRV32Config.fir@119722.4]
  assign cmd_read = _T_1829 | _T_1846; // @[Consts.scala 82:75:freechips.rocketchip.system.DefaultRV32Config.fir@119723.4]
  assign _T_1847 = io_req_bits_cmd == 5'h1; // @[Consts.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@119724.4]
  assign _T_1848 = io_req_bits_cmd == 5'h11; // @[Consts.scala 83:49:freechips.rocketchip.system.DefaultRV32Config.fir@119725.4]
  assign _T_1849 = _T_1847 | _T_1848; // @[Consts.scala 83:42:freechips.rocketchip.system.DefaultRV32Config.fir@119726.4]
  assign _T_1851 = _T_1849 | _T_1807; // @[Consts.scala 83:59:freechips.rocketchip.system.DefaultRV32Config.fir@119728.4]
  assign cmd_write = _T_1851 | _T_1846; // @[Consts.scala 83:76:freechips.rocketchip.system.DefaultRV32Config.fir@119746.4]
  assign _T_1869 = io_req_bits_cmd == 5'h5; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119747.4]
  assign _T_1870 = io_req_bits_cmd == 5'h17; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@119748.4]
  assign _T_1871 = _T_1869 | _T_1870; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119749.4]
  assign cmd_write_perms = cmd_write | _T_1871; // @[TLB.scala 285:35:freechips.rocketchip.system.DefaultRV32Config.fir@119750.4]
  assign _T_1872 = misaligned ? eff_array : 14'h0; // @[TLB.scala 290:8:freechips.rocketchip.system.DefaultRV32Config.fir@119752.4]
  assign _T_1873 = ~ c_array; // @[TLB.scala 291:19:freechips.rocketchip.system.DefaultRV32Config.fir@119753.4]
  assign _T_1874 = cmd_lrsc ? _T_1873 : 14'h0; // @[TLB.scala 291:8:freechips.rocketchip.system.DefaultRV32Config.fir@119754.4]
  assign ae_array = _T_1872 | _T_1874; // @[TLB.scala 290:37:freechips.rocketchip.system.DefaultRV32Config.fir@119755.4]
  assign _T_1875 = ~ pr_array; // @[TLB.scala 292:46:freechips.rocketchip.system.DefaultRV32Config.fir@119756.4]
  assign _T_1876 = ae_array | _T_1875; // @[TLB.scala 292:44:freechips.rocketchip.system.DefaultRV32Config.fir@119757.4]
  assign ae_ld_array = cmd_read ? _T_1876 : 14'h0; // @[TLB.scala 292:24:freechips.rocketchip.system.DefaultRV32Config.fir@119758.4]
  assign _T_1877 = ~ pw_array; // @[TLB.scala 294:37:freechips.rocketchip.system.DefaultRV32Config.fir@119759.4]
  assign _T_1878 = ae_array | _T_1877; // @[TLB.scala 294:35:freechips.rocketchip.system.DefaultRV32Config.fir@119760.4]
  assign _T_1879 = cmd_write_perms ? _T_1878 : 14'h0; // @[TLB.scala 294:8:freechips.rocketchip.system.DefaultRV32Config.fir@119761.4]
  assign _T_1880 = ~ pal_array_if_cached; // @[TLB.scala 295:26:freechips.rocketchip.system.DefaultRV32Config.fir@119762.4]
  assign _T_1881 = cmd_amo_logical ? _T_1880 : 14'h0; // @[TLB.scala 295:8:freechips.rocketchip.system.DefaultRV32Config.fir@119763.4]
  assign _T_1882 = _T_1879 | _T_1881; // @[TLB.scala 294:53:freechips.rocketchip.system.DefaultRV32Config.fir@119764.4]
  assign _T_1883 = ~ paa_array_if_cached; // @[TLB.scala 296:29:freechips.rocketchip.system.DefaultRV32Config.fir@119765.4]
  assign _T_1884 = cmd_amo_arithmetic ? _T_1883 : 14'h0; // @[TLB.scala 296:8:freechips.rocketchip.system.DefaultRV32Config.fir@119766.4]
  assign ae_st_array = _T_1882 | _T_1884; // @[TLB.scala 295:53:freechips.rocketchip.system.DefaultRV32Config.fir@119767.4]
  assign _T_1892 = misaligned & cmd_read; // @[TLB.scala 301:36:freechips.rocketchip.system.DefaultRV32Config.fir@119776.4]
  assign _T_1893 = ~ eff_array; // @[TLB.scala 301:49:freechips.rocketchip.system.DefaultRV32Config.fir@119777.4]
  assign ma_ld_array = _T_1892 ? _T_1893 : 14'h0; // @[TLB.scala 301:24:freechips.rocketchip.system.DefaultRV32Config.fir@119778.4]
  assign _T_1894 = misaligned & cmd_write; // @[TLB.scala 302:36:freechips.rocketchip.system.DefaultRV32Config.fir@119779.4]
  assign ma_st_array = _T_1894 ? _T_1893 : 14'h0; // @[TLB.scala 302:24:freechips.rocketchip.system.DefaultRV32Config.fir@119781.4]
  assign _T_1896 = r_array | ptw_ae_array; // @[TLB.scala 303:45:freechips.rocketchip.system.DefaultRV32Config.fir@119782.4]
  assign _T_1897 = ~ _T_1896; // @[TLB.scala 303:35:freechips.rocketchip.system.DefaultRV32Config.fir@119783.4]
  assign pf_ld_array = cmd_read ? _T_1897 : 14'h0; // @[TLB.scala 303:24:freechips.rocketchip.system.DefaultRV32Config.fir@119784.4]
  assign _T_1898 = w_array | ptw_ae_array; // @[TLB.scala 304:52:freechips.rocketchip.system.DefaultRV32Config.fir@119785.4]
  assign _T_1899 = ~ _T_1898; // @[TLB.scala 304:42:freechips.rocketchip.system.DefaultRV32Config.fir@119786.4]
  assign pf_st_array = cmd_write_perms ? _T_1899 : 14'h0; // @[TLB.scala 304:24:freechips.rocketchip.system.DefaultRV32Config.fir@119787.4]
  assign tlb_hit = real_hits != 13'h0; // @[TLB.scala 307:27:freechips.rocketchip.system.DefaultRV32Config.fir@119790.4]
  assign _T_1903 = tlb_hit == 1'h0; // @[TLB.scala 308:43:freechips.rocketchip.system.DefaultRV32Config.fir@119793.4]
  assign tlb_miss = vm_enabled & _T_1903; // @[TLB.scala 308:40:freechips.rocketchip.system.DefaultRV32Config.fir@119794.4]
  assign _T_1906 = io_req_valid & vm_enabled; // @[TLB.scala 312:22:freechips.rocketchip.system.DefaultRV32Config.fir@119797.4]
  assign _T_1907 = sector_hits_0 | sector_hits_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119799.6]
  assign _T_1908 = _T_1907 | sector_hits_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119800.6]
  assign _T_1909 = _T_1908 | sector_hits_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119801.6]
  assign _T_1910 = _T_1909 | sector_hits_4; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119802.6]
  assign _T_1911 = _T_1910 | sector_hits_5; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119803.6]
  assign _T_1912 = _T_1911 | sector_hits_6; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119804.6]
  assign _T_1913 = _T_1912 | sector_hits_7; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119805.6]
  assign _T_1920 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119813.8]
  assign _T_1921 = _T_1920[7:4]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@119814.8]
  assign _T_1922 = _T_1920[3:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@119815.8]
  assign _T_1923 = _T_1921 != 4'h0; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@119816.8]
  assign _T_1924 = _T_1921 | _T_1922; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@119817.8]
  assign _T_1925 = _T_1924[3:2]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@119818.8]
  assign _T_1926 = _T_1924[1:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@119819.8]
  assign _T_1927 = _T_1925 != 2'h0; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@119820.8]
  assign _T_1928 = _T_1925 | _T_1926; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@119821.8]
  assign _T_1929 = _T_1928[1]; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@119822.8]
  assign _T_1931 = {_T_1923,_T_1927,_T_1929}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119824.8]
  assign _T_1932 = {_T_1904, 1'h0}; // @[Replacement.scala 46:28:freechips.rocketchip.system.DefaultRV32Config.fir@119825.8]
  assign _T_1933 = _T_1931[2]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119826.8]
  assign _T_1934 = _T_1933 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119827.8]
  assign _T_1936 = _T_1932 | 8'h2; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119829.8]
  assign _T_1937 = ~ _T_1932; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119830.8]
  assign _T_1938 = _T_1937 | 8'h2; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119831.8]
  assign _T_1939 = ~ _T_1938; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119832.8]
  assign _T_1940 = _T_1934 ? _T_1936 : _T_1939; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119833.8]
  assign _T_1941 = {1'h1,_T_1933}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119834.8]
  assign _T_1942 = _T_1931[1]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119835.8]
  assign _T_1943 = _T_1942 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119836.8]
  assign _T_1944 = 4'h1 << _T_1941; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119837.8]
  assign _GEN_983 = {{4'd0}, _T_1944}; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119838.8]
  assign _T_1945 = _T_1940 | _GEN_983; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119838.8]
  assign _T_1946 = ~ _T_1940; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119839.8]
  assign _T_1947 = _T_1946 | _GEN_983; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119840.8]
  assign _T_1948 = ~ _T_1947; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119841.8]
  assign _T_1949 = _T_1943 ? _T_1945 : _T_1948; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119842.8]
  assign _T_1950 = {1'h1,_T_1933,_T_1942}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119843.8]
  assign _T_1951 = _T_1931[0]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119844.8]
  assign _T_1952 = _T_1951 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119845.8]
  assign _T_1953 = 8'h1 << _T_1950; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119846.8]
  assign _T_1954 = _T_1949 | _T_1953; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119847.8]
  assign _T_1955 = ~ _T_1949; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119848.8]
  assign _T_1956 = _T_1955 | _T_1953; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119849.8]
  assign _T_1957 = ~ _T_1956; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119850.8]
  assign _T_1958 = _T_1952 ? _T_1954 : _T_1957; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119851.8]
  assign _T_1960 = _T_1958[7:1]; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@119853.8]
  assign _T_1961 = superpage_hits_0 | superpage_hits_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119856.6]
  assign _T_1962 = _T_1961 | superpage_hits_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119857.6]
  assign _T_1963 = _T_1962 | superpage_hits_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@119858.6]
  assign _T_1966 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119862.8]
  assign _T_1967 = _T_1966[3:2]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@119863.8]
  assign _T_1968 = _T_1966[1:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@119864.8]
  assign _T_1969 = _T_1967 != 2'h0; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@119865.8]
  assign _T_1970 = _T_1967 | _T_1968; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@119866.8]
  assign _T_1971 = _T_1970[1]; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@119867.8]
  assign _T_1972 = {_T_1969,_T_1971}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119868.8]
  assign _T_1973 = {_T_1905, 1'h0}; // @[Replacement.scala 46:28:freechips.rocketchip.system.DefaultRV32Config.fir@119869.8]
  assign _T_1974 = _T_1972[1]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119870.8]
  assign _T_1975 = _T_1974 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119871.8]
  assign _T_1977 = _T_1973 | 4'h2; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119873.8]
  assign _T_1978 = ~ _T_1973; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119874.8]
  assign _T_1979 = _T_1978 | 4'h2; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119875.8]
  assign _T_1980 = ~ _T_1979; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119876.8]
  assign _T_1981 = _T_1975 ? _T_1977 : _T_1980; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119877.8]
  assign _T_1982 = {1'h1,_T_1974}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@119878.8]
  assign _T_1983 = _T_1972[0]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@119879.8]
  assign _T_1984 = _T_1983 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@119880.8]
  assign _T_1985 = 4'h1 << _T_1982; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119881.8]
  assign _T_1986 = _T_1981 | _T_1985; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119882.8]
  assign _T_1987 = ~ _T_1981; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119883.8]
  assign _T_1988 = _T_1987 | _T_1985; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119884.8]
  assign _T_1989 = ~ _T_1988; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119885.8]
  assign _T_1990 = _T_1984 ? _T_1986 : _T_1989; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@119886.8]
  assign _T_1992 = _T_1990[3:1]; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@119888.8]
  assign _T_1993 = real_hits[5:0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119892.4]
  assign _T_1994 = _T_1993[2:0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119893.4]
  assign _T_1995 = _T_1994[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119894.4]
  assign _T_1997 = _T_1994[2:1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119896.4]
  assign _T_1998 = _T_1997[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119897.4]
  assign _T_2000 = _T_1997[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119899.4]
  assign _T_2002 = _T_1998 | _T_2000; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119901.4]
  assign _T_2004 = _T_1998 & _T_2000; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119903.4]
  assign _T_2006 = _T_1995 | _T_2002; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119905.4]
  assign _T_2008 = _T_1995 & _T_2002; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119907.4]
  assign _T_2009 = _T_2004 | _T_2008; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119908.4]
  assign _T_2010 = _T_1993[5:3]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119909.4]
  assign _T_2011 = _T_2010[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119910.4]
  assign _T_2013 = _T_2010[2:1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119912.4]
  assign _T_2014 = _T_2013[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119913.4]
  assign _T_2016 = _T_2013[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119915.4]
  assign _T_2018 = _T_2014 | _T_2016; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119917.4]
  assign _T_2020 = _T_2014 & _T_2016; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119919.4]
  assign _T_2022 = _T_2011 | _T_2018; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119921.4]
  assign _T_2024 = _T_2011 & _T_2018; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119923.4]
  assign _T_2025 = _T_2020 | _T_2024; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119924.4]
  assign _T_2026 = _T_2006 | _T_2022; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119925.4]
  assign _T_2027 = _T_2009 | _T_2025; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@119926.4]
  assign _T_2028 = _T_2006 & _T_2022; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119927.4]
  assign _T_2029 = _T_2027 | _T_2028; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119928.4]
  assign _T_2030 = real_hits[12:6]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119929.4]
  assign _T_2031 = _T_2030[2:0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119930.4]
  assign _T_2032 = _T_2031[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119931.4]
  assign _T_2034 = _T_2031[2:1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119933.4]
  assign _T_2035 = _T_2034[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119934.4]
  assign _T_2037 = _T_2034[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119936.4]
  assign _T_2039 = _T_2035 | _T_2037; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119938.4]
  assign _T_2041 = _T_2035 & _T_2037; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119940.4]
  assign _T_2043 = _T_2032 | _T_2039; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119942.4]
  assign _T_2045 = _T_2032 & _T_2039; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119944.4]
  assign _T_2046 = _T_2041 | _T_2045; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119945.4]
  assign _T_2047 = _T_2030[6:3]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119946.4]
  assign _T_2048 = _T_2047[1:0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119947.4]
  assign _T_2049 = _T_2048[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119948.4]
  assign _T_2051 = _T_2048[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119950.4]
  assign _T_2053 = _T_2049 | _T_2051; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119952.4]
  assign _T_2055 = _T_2049 & _T_2051; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119954.4]
  assign _T_2057 = _T_2047[3:2]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119956.4]
  assign _T_2058 = _T_2057[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@119957.4]
  assign _T_2060 = _T_2057[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@119959.4]
  assign _T_2062 = _T_2058 | _T_2060; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119961.4]
  assign _T_2064 = _T_2058 & _T_2060; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119963.4]
  assign _T_2066 = _T_2053 | _T_2062; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119965.4]
  assign _T_2067 = _T_2055 | _T_2064; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@119966.4]
  assign _T_2068 = _T_2053 & _T_2062; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119967.4]
  assign _T_2069 = _T_2067 | _T_2068; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119968.4]
  assign _T_2070 = _T_2043 | _T_2066; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@119969.4]
  assign _T_2071 = _T_2046 | _T_2069; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@119970.4]
  assign _T_2072 = _T_2043 & _T_2066; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119971.4]
  assign _T_2073 = _T_2071 | _T_2072; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119972.4]
  assign _T_2075 = _T_2029 | _T_2073; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@119974.4]
  assign _T_2076 = _T_2026 & _T_2070; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@119975.4]
  assign multipleHits = _T_2075 | _T_2076; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@119976.4]
  assign _T_2079 = pf_ld_array & hits; // @[TLB.scala 325:57:freechips.rocketchip.system.DefaultRV32Config.fir@119980.4]
  assign _T_2083 = pf_st_array & hits; // @[TLB.scala 326:64:freechips.rocketchip.system.DefaultRV32Config.fir@119985.4]
  assign _T_2089 = ae_ld_array & hits; // @[TLB.scala 328:33:freechips.rocketchip.system.DefaultRV32Config.fir@119993.4]
  assign _T_2091 = ae_st_array & hits; // @[TLB.scala 329:33:freechips.rocketchip.system.DefaultRV32Config.fir@119996.4]
  assign _T_2096 = ma_ld_array & hits; // @[TLB.scala 331:33:freechips.rocketchip.system.DefaultRV32Config.fir@120003.4]
  assign _T_2098 = ma_st_array & hits; // @[TLB.scala 332:33:freechips.rocketchip.system.DefaultRV32Config.fir@120006.4]
  assign _T_2100 = c_array & hits; // @[TLB.scala 334:33:freechips.rocketchip.system.DefaultRV32Config.fir@120010.4]
  assign _T_2107 = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 337:29:freechips.rocketchip.system.DefaultRV32Config.fir@120020.4]
  assign _T_2113 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@120031.4]
  assign _T_2114 = _T_2113 & tlb_miss; // @[TLB.scala 346:25:freechips.rocketchip.system.DefaultRV32Config.fir@120032.4]
  assign _GEN_985 = _T_1973[3:1]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120040.6]
  assign _T_2119 = {{1'd0}, _GEN_985}; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120040.6]
  assign _T_2120 = _T_2119[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120041.6]
  assign _T_2122 = {1'h1,_T_2120}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120043.6]
  assign _T_2126 = _T_1973 >> _T_2122; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120047.6]
  assign _T_2127 = _T_2126[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120048.6]
  assign _T_2129 = {1'h1,_T_2120,_T_2127}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120050.6]
  assign _T_2130 = _T_2129[1:0]; // @[Replacement.scala 63:8:freechips.rocketchip.system.DefaultRV32Config.fir@120051.6]
  assign _T_2133 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120054.6]
  assign _T_2134 = _T_2133 == 4'hf; // @[TLB.scala 394:16:freechips.rocketchip.system.DefaultRV32Config.fir@120055.6]
  assign _T_2135 = ~ _T_2133; // @[TLB.scala 394:43:freechips.rocketchip.system.DefaultRV32Config.fir@120056.6]
  assign _T_2136 = _T_2135[0]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120057.6]
  assign _T_2137 = _T_2135[1]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120058.6]
  assign _T_2138 = _T_2135[2]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120059.6]
  assign _GEN_986 = _T_1932[7:1]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120070.6]
  assign _T_2148 = {{1'd0}, _GEN_986}; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120070.6]
  assign _T_2149 = _T_2148[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120071.6]
  assign _T_2151 = {1'h1,_T_2149}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120073.6]
  assign _T_2155 = _T_1932 >> _T_2151; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120077.6]
  assign _T_2156 = _T_2155[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120078.6]
  assign _T_2158 = {1'h1,_T_2149,_T_2156}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120080.6]
  assign _T_2162 = _T_1932 >> _T_2158; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120084.6]
  assign _T_2163 = _T_2162[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@120085.6]
  assign _T_2165 = {1'h1,_T_2149,_T_2156,_T_2163}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120087.6]
  assign _T_2166 = _T_2165[2:0]; // @[Replacement.scala 63:8:freechips.rocketchip.system.DefaultRV32Config.fir@120088.6]
  assign _T_2197 = {_T_421,_T_415,_T_409,_T_403,_T_397,_T_391,_T_385,_T_379}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@120119.6]
  assign _T_2198 = _T_2197 == 8'hff; // @[TLB.scala 394:16:freechips.rocketchip.system.DefaultRV32Config.fir@120120.6]
  assign _T_2199 = ~ _T_2197; // @[TLB.scala 394:43:freechips.rocketchip.system.DefaultRV32Config.fir@120121.6]
  assign _T_2200 = _T_2199[0]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120122.6]
  assign _T_2201 = _T_2199[1]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120123.6]
  assign _T_2202 = _T_2199[2]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120124.6]
  assign _T_2203 = _T_2199[3]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120125.6]
  assign _T_2204 = _T_2199[4]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120126.6]
  assign _T_2205 = _T_2199[5]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120127.6]
  assign _T_2206 = _T_2199[6]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@120128.6]
  assign _T_2243 = state == 2'h2; // @[TLB.scala 360:17:freechips.rocketchip.system.DefaultRV32Config.fir@120180.4]
  assign _T_2244 = _T_2243 & io_sfence_valid; // @[TLB.scala 360:28:freechips.rocketchip.system.DefaultRV32Config.fir@120181.4]
  assign _T_2245 = io_sfence_bits_rs1 == 1'h0; // @[TLB.scala 368:14:freechips.rocketchip.system.DefaultRV32Config.fir@120189.6]
  assign _T_2246 = io_sfence_bits_addr[31:12]; // @[TLB.scala 368:58:freechips.rocketchip.system.DefaultRV32Config.fir@120190.6]
  assign _T_2247 = _T_2246 == vpn; // @[TLB.scala 368:72:freechips.rocketchip.system.DefaultRV32Config.fir@120191.6]
  assign _T_2248 = _T_2245 | _T_2247; // @[TLB.scala 368:34:freechips.rocketchip.system.DefaultRV32Config.fir@120192.6]
  assign _T_2250 = _T_2248 | reset; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@120194.6]
  assign _T_2251 = _T_2250 == 1'h0; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@120195.6]
  assign _T_2257 = _T_380[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@120209.8]
  assign _T_2258 = _T_2257 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@120210.8]
  assign _T_2261 = sectored_entries_0_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120217.10]
  assign _T_2273 = sectored_entries_0_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120241.10]
  assign _T_2278 = sectored_entries_0_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120252.10]
  assign _T_2290 = sectored_entries_0_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120276.10]
  assign _T_2295 = sectored_entries_0_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120287.10]
  assign _T_2307 = sectored_entries_0_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120311.10]
  assign _T_2312 = sectored_entries_0_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120322.10]
  assign _T_2324 = sectored_entries_0_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120346.10]
  assign _T_2395 = _T_2273 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120508.10]
  assign _GEN_648 = _T_2395 ? 1'h0 : _GEN_472; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120509.10]
  assign _T_2396 = _T_2290 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120512.10]
  assign _GEN_649 = _T_2396 ? 1'h0 : _GEN_473; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120513.10]
  assign _T_2397 = _T_2307 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120516.10]
  assign _GEN_650 = _T_2397 ? 1'h0 : _GEN_474; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120517.10]
  assign _T_2398 = _T_2324 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120520.10]
  assign _GEN_651 = _T_2398 ? 1'h0 : _GEN_475; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120521.10]
  assign _GEN_652 = io_sfence_bits_rs2 & _GEN_648; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120367.8]
  assign _GEN_653 = io_sfence_bits_rs2 & _GEN_649; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120367.8]
  assign _GEN_654 = io_sfence_bits_rs2 & _GEN_650; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120367.8]
  assign _GEN_655 = io_sfence_bits_rs2 & _GEN_651; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120367.8]
  assign _T_2404 = _T_386[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@120540.8]
  assign _T_2405 = _T_2404 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@120541.8]
  assign _T_2408 = sectored_entries_1_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120548.10]
  assign _T_2420 = sectored_entries_1_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120572.10]
  assign _T_2425 = sectored_entries_1_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120583.10]
  assign _T_2437 = sectored_entries_1_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120607.10]
  assign _T_2442 = sectored_entries_1_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120618.10]
  assign _T_2454 = sectored_entries_1_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120642.10]
  assign _T_2459 = sectored_entries_1_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120653.10]
  assign _T_2471 = sectored_entries_1_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120677.10]
  assign _T_2542 = _T_2420 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120839.10]
  assign _GEN_676 = _T_2542 ? 1'h0 : _GEN_482; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120840.10]
  assign _T_2543 = _T_2437 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120843.10]
  assign _GEN_677 = _T_2543 ? 1'h0 : _GEN_483; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120844.10]
  assign _T_2544 = _T_2454 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120847.10]
  assign _GEN_678 = _T_2544 ? 1'h0 : _GEN_484; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120848.10]
  assign _T_2545 = _T_2471 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@120851.10]
  assign _GEN_679 = _T_2545 ? 1'h0 : _GEN_485; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@120852.10]
  assign _GEN_680 = io_sfence_bits_rs2 & _GEN_676; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120698.8]
  assign _GEN_681 = io_sfence_bits_rs2 & _GEN_677; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120698.8]
  assign _GEN_682 = io_sfence_bits_rs2 & _GEN_678; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120698.8]
  assign _GEN_683 = io_sfence_bits_rs2 & _GEN_679; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@120698.8]
  assign _T_2551 = _T_392[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@120871.8]
  assign _T_2552 = _T_2551 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@120872.8]
  assign _T_2555 = sectored_entries_2_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120879.10]
  assign _T_2567 = sectored_entries_2_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120903.10]
  assign _T_2572 = sectored_entries_2_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120914.10]
  assign _T_2584 = sectored_entries_2_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120938.10]
  assign _T_2589 = sectored_entries_2_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120949.10]
  assign _T_2601 = sectored_entries_2_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120973.10]
  assign _T_2606 = sectored_entries_2_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@120984.10]
  assign _T_2618 = sectored_entries_2_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121008.10]
  assign _T_2689 = _T_2567 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121170.10]
  assign _GEN_704 = _T_2689 ? 1'h0 : _GEN_492; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121171.10]
  assign _T_2690 = _T_2584 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121174.10]
  assign _GEN_705 = _T_2690 ? 1'h0 : _GEN_493; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121175.10]
  assign _T_2691 = _T_2601 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121178.10]
  assign _GEN_706 = _T_2691 ? 1'h0 : _GEN_494; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121179.10]
  assign _T_2692 = _T_2618 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121182.10]
  assign _GEN_707 = _T_2692 ? 1'h0 : _GEN_495; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121183.10]
  assign _GEN_708 = io_sfence_bits_rs2 & _GEN_704; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121029.8]
  assign _GEN_709 = io_sfence_bits_rs2 & _GEN_705; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121029.8]
  assign _GEN_710 = io_sfence_bits_rs2 & _GEN_706; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121029.8]
  assign _GEN_711 = io_sfence_bits_rs2 & _GEN_707; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121029.8]
  assign _T_2698 = _T_398[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@121202.8]
  assign _T_2699 = _T_2698 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@121203.8]
  assign _T_2702 = sectored_entries_3_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121210.10]
  assign _T_2714 = sectored_entries_3_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121234.10]
  assign _T_2719 = sectored_entries_3_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121245.10]
  assign _T_2731 = sectored_entries_3_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121269.10]
  assign _T_2736 = sectored_entries_3_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121280.10]
  assign _T_2748 = sectored_entries_3_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121304.10]
  assign _T_2753 = sectored_entries_3_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121315.10]
  assign _T_2765 = sectored_entries_3_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121339.10]
  assign _T_2836 = _T_2714 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121501.10]
  assign _GEN_732 = _T_2836 ? 1'h0 : _GEN_502; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121502.10]
  assign _T_2837 = _T_2731 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121505.10]
  assign _GEN_733 = _T_2837 ? 1'h0 : _GEN_503; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121506.10]
  assign _T_2838 = _T_2748 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121509.10]
  assign _GEN_734 = _T_2838 ? 1'h0 : _GEN_504; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121510.10]
  assign _T_2839 = _T_2765 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121513.10]
  assign _GEN_735 = _T_2839 ? 1'h0 : _GEN_505; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121514.10]
  assign _GEN_736 = io_sfence_bits_rs2 & _GEN_732; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121360.8]
  assign _GEN_737 = io_sfence_bits_rs2 & _GEN_733; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121360.8]
  assign _GEN_738 = io_sfence_bits_rs2 & _GEN_734; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121360.8]
  assign _GEN_739 = io_sfence_bits_rs2 & _GEN_735; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121360.8]
  assign _T_2845 = _T_404[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@121533.8]
  assign _T_2846 = _T_2845 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@121534.8]
  assign _T_2849 = sectored_entries_4_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121541.10]
  assign _T_2861 = sectored_entries_4_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121565.10]
  assign _T_2866 = sectored_entries_4_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121576.10]
  assign _T_2878 = sectored_entries_4_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121600.10]
  assign _T_2883 = sectored_entries_4_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121611.10]
  assign _T_2895 = sectored_entries_4_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121635.10]
  assign _T_2900 = sectored_entries_4_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121646.10]
  assign _T_2912 = sectored_entries_4_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121670.10]
  assign _T_2983 = _T_2861 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121832.10]
  assign _GEN_760 = _T_2983 ? 1'h0 : _GEN_512; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121833.10]
  assign _T_2984 = _T_2878 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121836.10]
  assign _GEN_761 = _T_2984 ? 1'h0 : _GEN_513; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121837.10]
  assign _T_2985 = _T_2895 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121840.10]
  assign _GEN_762 = _T_2985 ? 1'h0 : _GEN_514; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121841.10]
  assign _T_2986 = _T_2912 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@121844.10]
  assign _GEN_763 = _T_2986 ? 1'h0 : _GEN_515; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@121845.10]
  assign _GEN_764 = io_sfence_bits_rs2 & _GEN_760; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121691.8]
  assign _GEN_765 = io_sfence_bits_rs2 & _GEN_761; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121691.8]
  assign _GEN_766 = io_sfence_bits_rs2 & _GEN_762; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121691.8]
  assign _GEN_767 = io_sfence_bits_rs2 & _GEN_763; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@121691.8]
  assign _T_2992 = _T_410[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@121864.8]
  assign _T_2993 = _T_2992 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@121865.8]
  assign _T_2996 = sectored_entries_5_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121872.10]
  assign _T_3008 = sectored_entries_5_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121896.10]
  assign _T_3013 = sectored_entries_5_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121907.10]
  assign _T_3025 = sectored_entries_5_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121931.10]
  assign _T_3030 = sectored_entries_5_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121942.10]
  assign _T_3042 = sectored_entries_5_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121966.10]
  assign _T_3047 = sectored_entries_5_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@121977.10]
  assign _T_3059 = sectored_entries_5_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122001.10]
  assign _T_3130 = _T_3008 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122163.10]
  assign _GEN_788 = _T_3130 ? 1'h0 : _GEN_522; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122164.10]
  assign _T_3131 = _T_3025 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122167.10]
  assign _GEN_789 = _T_3131 ? 1'h0 : _GEN_523; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122168.10]
  assign _T_3132 = _T_3042 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122171.10]
  assign _GEN_790 = _T_3132 ? 1'h0 : _GEN_524; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122172.10]
  assign _T_3133 = _T_3059 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122175.10]
  assign _GEN_791 = _T_3133 ? 1'h0 : _GEN_525; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122176.10]
  assign _GEN_792 = io_sfence_bits_rs2 & _GEN_788; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122022.8]
  assign _GEN_793 = io_sfence_bits_rs2 & _GEN_789; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122022.8]
  assign _GEN_794 = io_sfence_bits_rs2 & _GEN_790; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122022.8]
  assign _GEN_795 = io_sfence_bits_rs2 & _GEN_791; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122022.8]
  assign _T_3139 = _T_416[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@122195.8]
  assign _T_3140 = _T_3139 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@122196.8]
  assign _T_3143 = sectored_entries_6_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122203.10]
  assign _T_3155 = sectored_entries_6_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122227.10]
  assign _T_3160 = sectored_entries_6_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122238.10]
  assign _T_3172 = sectored_entries_6_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122262.10]
  assign _T_3177 = sectored_entries_6_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122273.10]
  assign _T_3189 = sectored_entries_6_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122297.10]
  assign _T_3194 = sectored_entries_6_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122308.10]
  assign _T_3206 = sectored_entries_6_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122332.10]
  assign _T_3277 = _T_3155 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122494.10]
  assign _GEN_816 = _T_3277 ? 1'h0 : _GEN_532; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122495.10]
  assign _T_3278 = _T_3172 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122498.10]
  assign _GEN_817 = _T_3278 ? 1'h0 : _GEN_533; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122499.10]
  assign _T_3279 = _T_3189 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122502.10]
  assign _GEN_818 = _T_3279 ? 1'h0 : _GEN_534; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122503.10]
  assign _T_3280 = _T_3206 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122506.10]
  assign _GEN_819 = _T_3280 ? 1'h0 : _GEN_535; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122507.10]
  assign _GEN_820 = io_sfence_bits_rs2 & _GEN_816; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122353.8]
  assign _GEN_821 = io_sfence_bits_rs2 & _GEN_817; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122353.8]
  assign _GEN_822 = io_sfence_bits_rs2 & _GEN_818; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122353.8]
  assign _GEN_823 = io_sfence_bits_rs2 & _GEN_819; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122353.8]
  assign _T_3286 = _T_422[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@122526.8]
  assign _T_3287 = _T_3286 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@122527.8]
  assign _T_3290 = sectored_entries_7_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122534.10]
  assign _T_3302 = sectored_entries_7_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122558.10]
  assign _T_3307 = sectored_entries_7_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122569.10]
  assign _T_3319 = sectored_entries_7_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122593.10]
  assign _T_3324 = sectored_entries_7_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122604.10]
  assign _T_3336 = sectored_entries_7_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122628.10]
  assign _T_3341 = sectored_entries_7_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122639.10]
  assign _T_3353 = sectored_entries_7_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@122663.10]
  assign _T_3424 = _T_3302 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122825.10]
  assign _GEN_844 = _T_3424 ? 1'h0 : _GEN_542; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122826.10]
  assign _T_3425 = _T_3319 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122829.10]
  assign _GEN_845 = _T_3425 ? 1'h0 : _GEN_543; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122830.10]
  assign _T_3426 = _T_3336 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122833.10]
  assign _GEN_846 = _T_3426 ? 1'h0 : _GEN_544; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122834.10]
  assign _T_3427 = _T_3353 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122837.10]
  assign _GEN_847 = _T_3427 ? 1'h0 : _GEN_545; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122838.10]
  assign _GEN_848 = io_sfence_bits_rs2 & _GEN_844; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122684.8]
  assign _GEN_849 = io_sfence_bits_rs2 & _GEN_845; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122684.8]
  assign _GEN_850 = io_sfence_bits_rs2 & _GEN_846; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122684.8]
  assign _GEN_851 = io_sfence_bits_rs2 & _GEN_847; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122684.8]
  assign _T_3459 = _T_758 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122904.10]
  assign _GEN_857 = _T_3459 ? 1'h0 : _GEN_458; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122905.10]
  assign _GEN_858 = io_sfence_bits_rs2 & _GEN_857; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122868.8]
  assign _T_3491 = _T_782 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@122968.10]
  assign _GEN_861 = _T_3491 ? 1'h0 : _GEN_462; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@122969.10]
  assign _GEN_862 = io_sfence_bits_rs2 & _GEN_861; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122932.8]
  assign _T_3523 = _T_806 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@123032.10]
  assign _GEN_865 = _T_3523 ? 1'h0 : _GEN_466; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@123033.10]
  assign _GEN_866 = io_sfence_bits_rs2 & _GEN_865; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@122996.8]
  assign _T_3555 = _T_830 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@123096.10]
  assign _GEN_869 = _T_3555 ? 1'h0 : _GEN_470; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@123097.10]
  assign _GEN_870 = io_sfence_bits_rs2 & _GEN_869; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@123060.8]
  assign _T_3587 = _T_21 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@123160.10]
  assign _GEN_873 = _T_3587 ? 1'h0 : _GEN_454; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@123161.10]
  assign _GEN_874 = io_sfence_bits_rs2 & _GEN_873; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@123124.8]
  assign _T_3589 = multipleHits | reset; // @[TLB.scala 375:24:freechips.rocketchip.system.DefaultRV32Config.fir@123170.4]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 324:16:freechips.rocketchip.system.DefaultRV32Config.fir@119978.4]
  assign io_resp_miss = _T_2107 | multipleHits; // @[TLB.scala 337:16:freechips.rocketchip.system.DefaultRV32Config.fir@120022.4]
  assign io_resp_paddr = {ppn,_T_33}; // @[TLB.scala 338:17:freechips.rocketchip.system.DefaultRV32Config.fir@120025.4]
  assign io_resp_pf_ld = _T_2079 != 14'h0; // @[TLB.scala 325:17:freechips.rocketchip.system.DefaultRV32Config.fir@119983.4]
  assign io_resp_pf_st = _T_2083 != 14'h0; // @[TLB.scala 326:17:freechips.rocketchip.system.DefaultRV32Config.fir@119988.4]
  assign io_resp_ae_ld = _T_2089 != 14'h0; // @[TLB.scala 328:17:freechips.rocketchip.system.DefaultRV32Config.fir@119995.4]
  assign io_resp_ae_st = _T_2091 != 14'h0; // @[TLB.scala 329:17:freechips.rocketchip.system.DefaultRV32Config.fir@119998.4]
  assign io_resp_ma_ld = _T_2096 != 14'h0; // @[TLB.scala 331:17:freechips.rocketchip.system.DefaultRV32Config.fir@120005.4]
  assign io_resp_ma_st = _T_2098 != 14'h0; // @[TLB.scala 332:17:freechips.rocketchip.system.DefaultRV32Config.fir@120008.4]
  assign io_resp_cacheable = _T_2100 != 14'h0; // @[TLB.scala 334:21:freechips.rocketchip.system.DefaultRV32Config.fir@120012.4]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 340:20:freechips.rocketchip.system.DefaultRV32Config.fir@120027.4]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 342:29:freechips.rocketchip.system.DefaultRV32Config.fir@120030.4]
  assign _2_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign _2_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@116785.4]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@116816.4]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116808.4]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116808.4]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116808.4]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116808.4]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116808.4]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116808.4]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116808.4]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116809.4]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116809.4]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116809.4]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116809.4]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116809.4]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116809.4]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116809.4]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116810.4]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116810.4]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116810.4]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116810.4]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116810.4]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116810.4]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116810.4]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116811.4]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116811.4]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116811.4]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116811.4]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116811.4]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116811.4]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116811.4]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116812.4]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116812.4]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116812.4]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116812.4]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116812.4]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116812.4]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116812.4]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116813.4]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116813.4]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116813.4]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116813.4]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116813.4]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116813.4]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116813.4]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116814.4]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116814.4]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116814.4]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116814.4]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116814.4]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116814.4]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116814.4]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116815.4]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116815.4]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116815.4]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116815.4]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116815.4]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116815.4]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@116815.4]
  assign pmp_io_addr = {mpu_ppn,_T_33}; // @[TLB.scala 190:15:freechips.rocketchip.system.DefaultRV32Config.fir@116806.4]
  assign _2_1_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_u = _GEN_35[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_px = _GEN_35[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_1_io_x_c = _GEN_35[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117471.4]
  assign _2_2_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_u = _GEN_39[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_px = _GEN_39[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_2_io_x_c = _GEN_39[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117512.4]
  assign _2_3_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_u = _GEN_43[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_px = _GEN_43[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_3_io_x_c = _GEN_43[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117553.4]
  assign _2_4_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_u = _GEN_47[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_px = _GEN_47[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_4_io_x_c = _GEN_47[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117594.4]
  assign _2_5_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_u = _GEN_51[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_px = _GEN_51[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_5_io_x_c = _GEN_51[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117635.4]
  assign _2_6_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_u = _GEN_55[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_px = _GEN_55[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_6_io_x_c = _GEN_55[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117676.4]
  assign _2_7_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_u = _GEN_59[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_px = _GEN_59[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_7_io_x_c = _GEN_59[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117717.4]
  assign _2_8_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_u = _GEN_63[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_px = _GEN_63[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_8_io_x_c = _GEN_63[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117758.4]
  assign _2_9_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_9_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117798.4]
  assign _2_10_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_10_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117845.4]
  assign _2_11_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_11_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117892.4]
  assign _2_12_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_12_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117939.4]
  assign _2_13_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_13_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@117986.4]
  assign _2_14_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_u = _GEN_35[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_px = _GEN_35[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_14_io_x_c = _GEN_35[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118451.4]
  assign _2_15_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_u = _GEN_39[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_px = _GEN_39[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_15_io_x_c = _GEN_39[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118492.4]
  assign _2_16_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_u = _GEN_43[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_px = _GEN_43[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_16_io_x_c = _GEN_43[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118533.4]
  assign _2_17_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_u = _GEN_47[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_px = _GEN_47[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_17_io_x_c = _GEN_47[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118574.4]
  assign _2_18_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_u = _GEN_51[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_px = _GEN_51[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_18_io_x_c = _GEN_51[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118615.4]
  assign _2_19_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_u = _GEN_55[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_px = _GEN_55[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_19_io_x_c = _GEN_55[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118656.4]
  assign _2_20_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_u = _GEN_59[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_px = _GEN_59[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_20_io_x_c = _GEN_59[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118697.4]
  assign _2_21_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_u = _GEN_63[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_px = _GEN_63[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_21_io_x_c = _GEN_63[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118738.4]
  assign _2_22_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_22_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118778.4]
  assign _2_23_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_23_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118818.4]
  assign _2_24_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_24_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118858.4]
  assign _2_25_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_25_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118898.4]
  assign _2_26_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_26_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118938.4]
  assign _2_27_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_u = _GEN_35[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_px = _GEN_35[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_27_io_x_c = _GEN_35[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@118979.4]
  assign _2_28_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_u = _GEN_39[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_px = _GEN_39[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_28_io_x_c = _GEN_39[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119020.4]
  assign _2_29_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_u = _GEN_43[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_px = _GEN_43[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_29_io_x_c = _GEN_43[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119061.4]
  assign _2_30_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_u = _GEN_47[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_px = _GEN_47[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_30_io_x_c = _GEN_47[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119102.4]
  assign _2_31_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_u = _GEN_51[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_px = _GEN_51[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_31_io_x_c = _GEN_51[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119143.4]
  assign _2_32_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_u = _GEN_55[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_px = _GEN_55[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_32_io_x_c = _GEN_55[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119184.4]
  assign _2_33_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_u = _GEN_59[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_px = _GEN_59[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_33_io_x_c = _GEN_59[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119225.4]
  assign _2_34_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_u = _GEN_63[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_px = _GEN_63[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_34_io_x_c = _GEN_63[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119266.4]
  assign _2_35_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_35_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119306.4]
  assign _2_36_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_36_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119346.4]
  assign _2_37_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_37_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119386.4]
  assign _2_38_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
  assign _2_38_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@119426.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_72[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_73[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_75[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_76[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_78[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_79[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_81[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_82[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  special_entry_level = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  special_entry_tag = _RAND_85[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_86[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  state = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  r_refill_tag = _RAND_89[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_90[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_92[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_sectored_hit = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1904 = _RAND_94[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1905 = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            sectored_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            if (2'h0 == _T_996) begin
              sectored_entries_0_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            if (2'h1 == _T_996) begin
              sectored_entries_0_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            if (2'h2 == _T_996) begin
              sectored_entries_0_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            if (2'h3 == _T_996) begin
              sectored_entries_0_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2258) begin
            if (_T_2261) begin
              sectored_entries_0_valid_0 <= 1'h0;
            end else begin
              if (_T_382) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_0_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_994) begin
                          sectored_entries_0_valid_0 <= _GEN_84;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_0 <= _GEN_84;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_382) begin
              if (2'h0 == _T_477) begin
                sectored_entries_0_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_0 <= _GEN_84;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_994) begin
                      sectored_entries_0_valid_0 <= _GEN_84;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_0_valid_0 <= _GEN_652;
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_472;
      end
    end
    if (_T_3589) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2258) begin
            if (_T_2278) begin
              sectored_entries_0_valid_1 <= 1'h0;
            end else begin
              if (_T_382) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_0_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_994) begin
                          sectored_entries_0_valid_1 <= _GEN_85;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_1 <= _GEN_85;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_382) begin
              if (2'h1 == _T_477) begin
                sectored_entries_0_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_1 <= _GEN_85;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_994) begin
                      sectored_entries_0_valid_1 <= _GEN_85;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_0_valid_1 <= _GEN_653;
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_473;
      end
    end
    if (_T_3589) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2258) begin
            if (_T_2295) begin
              sectored_entries_0_valid_2 <= 1'h0;
            end else begin
              if (_T_382) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_0_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_994) begin
                          sectored_entries_0_valid_2 <= _GEN_86;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_2 <= _GEN_86;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_382) begin
              if (2'h2 == _T_477) begin
                sectored_entries_0_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_2 <= _GEN_86;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_994) begin
                      sectored_entries_0_valid_2 <= _GEN_86;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_0_valid_2 <= _GEN_654;
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_474;
      end
    end
    if (_T_3589) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2258) begin
            if (_T_2312) begin
              sectored_entries_0_valid_3 <= 1'h0;
            end else begin
              if (_T_382) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_0_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_994) begin
                          sectored_entries_0_valid_3 <= _GEN_87;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_3 <= _GEN_87;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_382) begin
              if (2'h3 == _T_477) begin
                sectored_entries_0_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_3 <= _GEN_87;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_994) begin
                      sectored_entries_0_valid_3 <= _GEN_87;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_0_valid_3 <= _GEN_655;
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_475;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            sectored_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            if (2'h0 == _T_996) begin
              sectored_entries_1_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            if (2'h1 == _T_996) begin
              sectored_entries_1_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            if (2'h2 == _T_996) begin
              sectored_entries_1_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            if (2'h3 == _T_996) begin
              sectored_entries_1_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2405) begin
            if (_T_2408) begin
              sectored_entries_1_valid_0 <= 1'h0;
            end else begin
              if (_T_388) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_1_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1011) begin
                          sectored_entries_1_valid_0 <= _GEN_106;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_0 <= _GEN_106;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_388) begin
              if (2'h0 == _T_477) begin
                sectored_entries_1_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_0 <= _GEN_106;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1011) begin
                      sectored_entries_1_valid_0 <= _GEN_106;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_1_valid_0 <= _GEN_680;
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_482;
      end
    end
    if (_T_3589) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2405) begin
            if (_T_2425) begin
              sectored_entries_1_valid_1 <= 1'h0;
            end else begin
              if (_T_388) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_1_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1011) begin
                          sectored_entries_1_valid_1 <= _GEN_107;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_1 <= _GEN_107;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_388) begin
              if (2'h1 == _T_477) begin
                sectored_entries_1_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_1 <= _GEN_107;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1011) begin
                      sectored_entries_1_valid_1 <= _GEN_107;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_1_valid_1 <= _GEN_681;
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_483;
      end
    end
    if (_T_3589) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2405) begin
            if (_T_2442) begin
              sectored_entries_1_valid_2 <= 1'h0;
            end else begin
              if (_T_388) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_1_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1011) begin
                          sectored_entries_1_valid_2 <= _GEN_108;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_2 <= _GEN_108;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_388) begin
              if (2'h2 == _T_477) begin
                sectored_entries_1_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_2 <= _GEN_108;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1011) begin
                      sectored_entries_1_valid_2 <= _GEN_108;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_1_valid_2 <= _GEN_682;
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_484;
      end
    end
    if (_T_3589) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2405) begin
            if (_T_2459) begin
              sectored_entries_1_valid_3 <= 1'h0;
            end else begin
              if (_T_388) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_1_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1011) begin
                          sectored_entries_1_valid_3 <= _GEN_109;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_3 <= _GEN_109;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_388) begin
              if (2'h3 == _T_477) begin
                sectored_entries_1_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_3 <= _GEN_109;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1011) begin
                      sectored_entries_1_valid_3 <= _GEN_109;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_1_valid_3 <= _GEN_683;
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_485;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            sectored_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            if (2'h0 == _T_996) begin
              sectored_entries_2_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            if (2'h1 == _T_996) begin
              sectored_entries_2_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            if (2'h2 == _T_996) begin
              sectored_entries_2_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            if (2'h3 == _T_996) begin
              sectored_entries_2_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2552) begin
            if (_T_2555) begin
              sectored_entries_2_valid_0 <= 1'h0;
            end else begin
              if (_T_394) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_2_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1028) begin
                          sectored_entries_2_valid_0 <= _GEN_128;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_0 <= _GEN_128;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_394) begin
              if (2'h0 == _T_477) begin
                sectored_entries_2_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_0 <= _GEN_128;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1028) begin
                      sectored_entries_2_valid_0 <= _GEN_128;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_2_valid_0 <= _GEN_708;
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_492;
      end
    end
    if (_T_3589) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2552) begin
            if (_T_2572) begin
              sectored_entries_2_valid_1 <= 1'h0;
            end else begin
              if (_T_394) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_2_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1028) begin
                          sectored_entries_2_valid_1 <= _GEN_129;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_1 <= _GEN_129;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_394) begin
              if (2'h1 == _T_477) begin
                sectored_entries_2_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_1 <= _GEN_129;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1028) begin
                      sectored_entries_2_valid_1 <= _GEN_129;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_2_valid_1 <= _GEN_709;
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_493;
      end
    end
    if (_T_3589) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2552) begin
            if (_T_2589) begin
              sectored_entries_2_valid_2 <= 1'h0;
            end else begin
              if (_T_394) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_2_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1028) begin
                          sectored_entries_2_valid_2 <= _GEN_130;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_2 <= _GEN_130;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_394) begin
              if (2'h2 == _T_477) begin
                sectored_entries_2_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_2 <= _GEN_130;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1028) begin
                      sectored_entries_2_valid_2 <= _GEN_130;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_2_valid_2 <= _GEN_710;
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_494;
      end
    end
    if (_T_3589) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2552) begin
            if (_T_2606) begin
              sectored_entries_2_valid_3 <= 1'h0;
            end else begin
              if (_T_394) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_2_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1028) begin
                          sectored_entries_2_valid_3 <= _GEN_131;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_3 <= _GEN_131;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_394) begin
              if (2'h3 == _T_477) begin
                sectored_entries_2_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_3 <= _GEN_131;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1028) begin
                      sectored_entries_2_valid_3 <= _GEN_131;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_2_valid_3 <= _GEN_711;
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_495;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            sectored_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            if (2'h0 == _T_996) begin
              sectored_entries_3_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            if (2'h1 == _T_996) begin
              sectored_entries_3_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            if (2'h2 == _T_996) begin
              sectored_entries_3_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            if (2'h3 == _T_996) begin
              sectored_entries_3_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2699) begin
            if (_T_2702) begin
              sectored_entries_3_valid_0 <= 1'h0;
            end else begin
              if (_T_400) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_3_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1045) begin
                          sectored_entries_3_valid_0 <= _GEN_150;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_0 <= _GEN_150;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_400) begin
              if (2'h0 == _T_477) begin
                sectored_entries_3_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_0 <= _GEN_150;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1045) begin
                      sectored_entries_3_valid_0 <= _GEN_150;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_3_valid_0 <= _GEN_736;
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_502;
      end
    end
    if (_T_3589) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2699) begin
            if (_T_2719) begin
              sectored_entries_3_valid_1 <= 1'h0;
            end else begin
              if (_T_400) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_3_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1045) begin
                          sectored_entries_3_valid_1 <= _GEN_151;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_1 <= _GEN_151;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_400) begin
              if (2'h1 == _T_477) begin
                sectored_entries_3_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_1 <= _GEN_151;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1045) begin
                      sectored_entries_3_valid_1 <= _GEN_151;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_3_valid_1 <= _GEN_737;
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_503;
      end
    end
    if (_T_3589) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2699) begin
            if (_T_2736) begin
              sectored_entries_3_valid_2 <= 1'h0;
            end else begin
              if (_T_400) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_3_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1045) begin
                          sectored_entries_3_valid_2 <= _GEN_152;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_2 <= _GEN_152;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_400) begin
              if (2'h2 == _T_477) begin
                sectored_entries_3_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_2 <= _GEN_152;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1045) begin
                      sectored_entries_3_valid_2 <= _GEN_152;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_3_valid_2 <= _GEN_738;
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_504;
      end
    end
    if (_T_3589) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2699) begin
            if (_T_2753) begin
              sectored_entries_3_valid_3 <= 1'h0;
            end else begin
              if (_T_400) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_3_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1045) begin
                          sectored_entries_3_valid_3 <= _GEN_153;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_3 <= _GEN_153;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_400) begin
              if (2'h3 == _T_477) begin
                sectored_entries_3_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_3 <= _GEN_153;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1045) begin
                      sectored_entries_3_valid_3 <= _GEN_153;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_3_valid_3 <= _GEN_739;
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_505;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            sectored_entries_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            if (2'h0 == _T_996) begin
              sectored_entries_4_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            if (2'h1 == _T_996) begin
              sectored_entries_4_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            if (2'h2 == _T_996) begin
              sectored_entries_4_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            if (2'h3 == _T_996) begin
              sectored_entries_4_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2846) begin
            if (_T_2849) begin
              sectored_entries_4_valid_0 <= 1'h0;
            end else begin
              if (_T_406) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_4_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1062) begin
                          sectored_entries_4_valid_0 <= _GEN_172;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_0 <= _GEN_172;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_406) begin
              if (2'h0 == _T_477) begin
                sectored_entries_4_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_0 <= _GEN_172;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1062) begin
                      sectored_entries_4_valid_0 <= _GEN_172;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_4_valid_0 <= _GEN_764;
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_512;
      end
    end
    if (_T_3589) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2846) begin
            if (_T_2866) begin
              sectored_entries_4_valid_1 <= 1'h0;
            end else begin
              if (_T_406) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_4_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1062) begin
                          sectored_entries_4_valid_1 <= _GEN_173;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_1 <= _GEN_173;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_406) begin
              if (2'h1 == _T_477) begin
                sectored_entries_4_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_1 <= _GEN_173;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1062) begin
                      sectored_entries_4_valid_1 <= _GEN_173;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_4_valid_1 <= _GEN_765;
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_513;
      end
    end
    if (_T_3589) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2846) begin
            if (_T_2883) begin
              sectored_entries_4_valid_2 <= 1'h0;
            end else begin
              if (_T_406) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_4_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1062) begin
                          sectored_entries_4_valid_2 <= _GEN_174;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_2 <= _GEN_174;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_406) begin
              if (2'h2 == _T_477) begin
                sectored_entries_4_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_2 <= _GEN_174;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1062) begin
                      sectored_entries_4_valid_2 <= _GEN_174;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_4_valid_2 <= _GEN_766;
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_514;
      end
    end
    if (_T_3589) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2846) begin
            if (_T_2900) begin
              sectored_entries_4_valid_3 <= 1'h0;
            end else begin
              if (_T_406) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_4_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1062) begin
                          sectored_entries_4_valid_3 <= _GEN_175;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_3 <= _GEN_175;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_406) begin
              if (2'h3 == _T_477) begin
                sectored_entries_4_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_3 <= _GEN_175;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1062) begin
                      sectored_entries_4_valid_3 <= _GEN_175;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_4_valid_3 <= _GEN_767;
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_515;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            sectored_entries_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            if (2'h0 == _T_996) begin
              sectored_entries_5_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            if (2'h1 == _T_996) begin
              sectored_entries_5_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            if (2'h2 == _T_996) begin
              sectored_entries_5_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            if (2'h3 == _T_996) begin
              sectored_entries_5_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2993) begin
            if (_T_2996) begin
              sectored_entries_5_valid_0 <= 1'h0;
            end else begin
              if (_T_412) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_5_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1079) begin
                          sectored_entries_5_valid_0 <= _GEN_194;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_0 <= _GEN_194;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_412) begin
              if (2'h0 == _T_477) begin
                sectored_entries_5_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_0 <= _GEN_194;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1079) begin
                      sectored_entries_5_valid_0 <= _GEN_194;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_5_valid_0 <= _GEN_792;
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_522;
      end
    end
    if (_T_3589) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2993) begin
            if (_T_3013) begin
              sectored_entries_5_valid_1 <= 1'h0;
            end else begin
              if (_T_412) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_5_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1079) begin
                          sectored_entries_5_valid_1 <= _GEN_195;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_1 <= _GEN_195;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_412) begin
              if (2'h1 == _T_477) begin
                sectored_entries_5_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_1 <= _GEN_195;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1079) begin
                      sectored_entries_5_valid_1 <= _GEN_195;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_5_valid_1 <= _GEN_793;
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_523;
      end
    end
    if (_T_3589) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2993) begin
            if (_T_3030) begin
              sectored_entries_5_valid_2 <= 1'h0;
            end else begin
              if (_T_412) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_5_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1079) begin
                          sectored_entries_5_valid_2 <= _GEN_196;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_2 <= _GEN_196;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_412) begin
              if (2'h2 == _T_477) begin
                sectored_entries_5_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_2 <= _GEN_196;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1079) begin
                      sectored_entries_5_valid_2 <= _GEN_196;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_5_valid_2 <= _GEN_794;
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_524;
      end
    end
    if (_T_3589) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2993) begin
            if (_T_3047) begin
              sectored_entries_5_valid_3 <= 1'h0;
            end else begin
              if (_T_412) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_5_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1079) begin
                          sectored_entries_5_valid_3 <= _GEN_197;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_3 <= _GEN_197;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_412) begin
              if (2'h3 == _T_477) begin
                sectored_entries_5_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_3 <= _GEN_197;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1079) begin
                      sectored_entries_5_valid_3 <= _GEN_197;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_5_valid_3 <= _GEN_795;
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_525;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            sectored_entries_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            if (2'h0 == _T_996) begin
              sectored_entries_6_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            if (2'h1 == _T_996) begin
              sectored_entries_6_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            if (2'h2 == _T_996) begin
              sectored_entries_6_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            if (2'h3 == _T_996) begin
              sectored_entries_6_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3140) begin
            if (_T_3143) begin
              sectored_entries_6_valid_0 <= 1'h0;
            end else begin
              if (_T_418) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_6_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1096) begin
                          sectored_entries_6_valid_0 <= _GEN_216;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_0 <= _GEN_216;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_418) begin
              if (2'h0 == _T_477) begin
                sectored_entries_6_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_0 <= _GEN_216;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1096) begin
                      sectored_entries_6_valid_0 <= _GEN_216;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_6_valid_0 <= _GEN_820;
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_532;
      end
    end
    if (_T_3589) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3140) begin
            if (_T_3160) begin
              sectored_entries_6_valid_1 <= 1'h0;
            end else begin
              if (_T_418) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_6_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1096) begin
                          sectored_entries_6_valid_1 <= _GEN_217;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_1 <= _GEN_217;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_418) begin
              if (2'h1 == _T_477) begin
                sectored_entries_6_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_1 <= _GEN_217;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1096) begin
                      sectored_entries_6_valid_1 <= _GEN_217;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_6_valid_1 <= _GEN_821;
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_533;
      end
    end
    if (_T_3589) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3140) begin
            if (_T_3177) begin
              sectored_entries_6_valid_2 <= 1'h0;
            end else begin
              if (_T_418) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_6_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1096) begin
                          sectored_entries_6_valid_2 <= _GEN_218;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_2 <= _GEN_218;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_418) begin
              if (2'h2 == _T_477) begin
                sectored_entries_6_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_2 <= _GEN_218;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1096) begin
                      sectored_entries_6_valid_2 <= _GEN_218;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_6_valid_2 <= _GEN_822;
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_534;
      end
    end
    if (_T_3589) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3140) begin
            if (_T_3194) begin
              sectored_entries_6_valid_3 <= 1'h0;
            end else begin
              if (_T_418) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_6_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1096) begin
                          sectored_entries_6_valid_3 <= _GEN_219;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_3 <= _GEN_219;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_418) begin
              if (2'h3 == _T_477) begin
                sectored_entries_6_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_3 <= _GEN_219;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1096) begin
                      sectored_entries_6_valid_3 <= _GEN_219;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_6_valid_3 <= _GEN_823;
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_535;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            sectored_entries_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            if (2'h0 == _T_996) begin
              sectored_entries_7_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            if (2'h1 == _T_996) begin
              sectored_entries_7_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            if (2'h2 == _T_996) begin
              sectored_entries_7_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            if (2'h3 == _T_996) begin
              sectored_entries_7_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3287) begin
            if (_T_3290) begin
              sectored_entries_7_valid_0 <= 1'h0;
            end else begin
              if (_T_424) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_7_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1113) begin
                          sectored_entries_7_valid_0 <= _GEN_238;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_0 <= _GEN_238;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_424) begin
              if (2'h0 == _T_477) begin
                sectored_entries_7_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_0 <= _GEN_238;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1113) begin
                      sectored_entries_7_valid_0 <= _GEN_238;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_7_valid_0 <= _GEN_848;
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_542;
      end
    end
    if (_T_3589) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3287) begin
            if (_T_3307) begin
              sectored_entries_7_valid_1 <= 1'h0;
            end else begin
              if (_T_424) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_7_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1113) begin
                          sectored_entries_7_valid_1 <= _GEN_239;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_1 <= _GEN_239;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_424) begin
              if (2'h1 == _T_477) begin
                sectored_entries_7_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_1 <= _GEN_239;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1113) begin
                      sectored_entries_7_valid_1 <= _GEN_239;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_7_valid_1 <= _GEN_849;
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_543;
      end
    end
    if (_T_3589) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3287) begin
            if (_T_3324) begin
              sectored_entries_7_valid_2 <= 1'h0;
            end else begin
              if (_T_424) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_7_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1113) begin
                          sectored_entries_7_valid_2 <= _GEN_240;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_2 <= _GEN_240;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_424) begin
              if (2'h2 == _T_477) begin
                sectored_entries_7_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_2 <= _GEN_240;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1113) begin
                      sectored_entries_7_valid_2 <= _GEN_240;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_7_valid_2 <= _GEN_850;
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_544;
      end
    end
    if (_T_3589) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3287) begin
            if (_T_3341) begin
              sectored_entries_7_valid_3 <= 1'h0;
            end else begin
              if (_T_424) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_7_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1113) begin
                          sectored_entries_7_valid_3 <= _GEN_241;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_3 <= _GEN_241;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_424) begin
              if (2'h3 == _T_477) begin
                sectored_entries_7_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_3 <= _GEN_241;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1113) begin
                      sectored_entries_7_valid_3 <= _GEN_241;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_7_valid_3 <= _GEN_851;
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_545;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_933) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_933) begin
            superpage_entries_0_data_0 <= _T_931;
          end
        end
      end
    end
    if (_T_3589) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (superpage_hits_0) begin
            superpage_entries_0_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              if (!(_T_915)) begin
                if (_T_932) begin
                  superpage_entries_0_valid_0 <= _GEN_66;
                end
              end
            end
          end
        end else begin
          superpage_entries_0_valid_0 <= _GEN_858;
        end
      end else begin
        if (_T_893) begin
          if (!(_T_915)) begin
            if (_T_932) begin
              superpage_entries_0_valid_0 <= _GEN_66;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_948) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_948) begin
            superpage_entries_1_data_0 <= _T_931;
          end
        end
      end
    end
    if (_T_3589) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (superpage_hits_1) begin
            superpage_entries_1_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              if (!(_T_915)) begin
                if (_T_932) begin
                  superpage_entries_1_valid_0 <= _GEN_70;
                end
              end
            end
          end
        end else begin
          superpage_entries_1_valid_0 <= _GEN_862;
        end
      end else begin
        if (_T_893) begin
          if (!(_T_915)) begin
            if (_T_932) begin
              superpage_entries_1_valid_0 <= _GEN_70;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_963) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_963) begin
            superpage_entries_2_data_0 <= _T_931;
          end
        end
      end
    end
    if (_T_3589) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (superpage_hits_2) begin
            superpage_entries_2_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              if (!(_T_915)) begin
                if (_T_932) begin
                  superpage_entries_2_valid_0 <= _GEN_74;
                end
              end
            end
          end
        end else begin
          superpage_entries_2_valid_0 <= _GEN_866;
        end
      end else begin
        if (_T_893) begin
          if (!(_T_915)) begin
            if (_T_932) begin
              superpage_entries_2_valid_0 <= _GEN_74;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_978) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_978) begin
            superpage_entries_3_data_0 <= _T_931;
          end
        end
      end
    end
    if (_T_3589) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (superpage_hits_3) begin
            superpage_entries_3_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              if (!(_T_915)) begin
                if (_T_932) begin
                  superpage_entries_3_valid_0 <= _GEN_78;
                end
              end
            end
          end
        end else begin
          superpage_entries_3_valid_0 <= _GEN_870;
        end
      end else begin
        if (_T_893) begin
          if (!(_T_915)) begin
            if (_T_932) begin
              superpage_entries_3_valid_0 <= _GEN_78;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (_T_915) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (_T_893) begin
      if (_T_915) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (_T_893) begin
      if (_T_915) begin
        special_entry_data_0 <= _T_931;
      end
    end
    if (_T_3589) begin
      special_entry_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_586) begin
            special_entry_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              special_entry_valid_0 <= _GEN_354;
            end
          end
        end else begin
          special_entry_valid_0 <= _GEN_874;
        end
      end else begin
        if (_T_893) begin
          special_entry_valid_0 <= _GEN_354;
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (io_ptw_resp_valid) begin
        state <= 2'h0;
      end else begin
        if (_T_2244) begin
          state <= 2'h3;
        end else begin
          if (_T_4) begin
            if (io_ptw_req_ready) begin
              if (io_sfence_valid) begin
                state <= 2'h3;
              end else begin
                state <= 2'h2;
              end
            end else begin
              if (io_sfence_valid) begin
                state <= 2'h0;
              end else begin
                if (_T_2114) begin
                  state <= 2'h1;
                end
              end
            end
          end else begin
            if (_T_2114) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if (_T_2114) begin
      r_refill_tag <= vpn;
    end
    if (_T_2114) begin
      if (_T_2134) begin
        r_superpage_repl_addr <= _T_2130;
      end else begin
        if (_T_2136) begin
          r_superpage_repl_addr <= 2'h0;
        end else begin
          if (_T_2137) begin
            r_superpage_repl_addr <= 2'h1;
          end else begin
            if (_T_2138) begin
              r_superpage_repl_addr <= 2'h2;
            end else begin
              r_superpage_repl_addr <= 2'h3;
            end
          end
        end
      end
    end
    if (_T_2114) begin
      if (_T_2198) begin
        r_sectored_repl_addr <= _T_2166;
      end else begin
        if (_T_2200) begin
          r_sectored_repl_addr <= 3'h0;
        end else begin
          if (_T_2201) begin
            r_sectored_repl_addr <= 3'h1;
          end else begin
            if (_T_2202) begin
              r_sectored_repl_addr <= 3'h2;
            end else begin
              if (_T_2203) begin
                r_sectored_repl_addr <= 3'h3;
              end else begin
                if (_T_2204) begin
                  r_sectored_repl_addr <= 3'h4;
                end else begin
                  if (_T_2205) begin
                    r_sectored_repl_addr <= 3'h5;
                  end else begin
                    if (_T_2206) begin
                      r_sectored_repl_addr <= 3'h6;
                    end else begin
                      r_sectored_repl_addr <= 3'h7;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_2114) begin
      r_sectored_hit_addr <= _T_1931;
    end
    if (_T_2114) begin
      r_sectored_hit <= _T_1913;
    end
    if (_T_1906) begin
      if (_T_1913) begin
        _T_1904 <= _T_1960;
      end
    end
    if (_T_1906) begin
      if (_T_1963) begin
        _T_1905 <= _T_1992;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & _T_2251) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:368 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@120197.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & _T_2251) begin
          $fatal; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@120198.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
`endif // __TLB

