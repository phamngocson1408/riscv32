`include "include_module.v"
`ifdef ___3
module _3( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115485.2]
  input         io_in_0_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [11:0] io_in_0_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input         io_in_0_bits_write, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [31:0] io_in_0_bits_wdata, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [3:0]  io_in_0_bits_eccMask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [3:0]  io_in_0_bits_way_en, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output        io_in_1_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input         io_in_1_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [11:0] io_in_1_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input         io_in_1_bits_write, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [31:0] io_in_1_bits_wdata, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [3:0]  io_in_1_bits_eccMask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [3:0]  io_in_1_bits_way_en, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output        io_in_2_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input         io_in_2_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [11:0] io_in_2_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [31:0] io_in_2_bits_wdata, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [3:0]  io_in_2_bits_eccMask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output        io_in_3_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input         io_in_3_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [11:0] io_in_3_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [31:0] io_in_3_bits_wdata, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  input  [3:0]  io_in_3_bits_eccMask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output        io_out_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output [11:0] io_out_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output        io_out_bits_write, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output [31:0] io_out_bits_wdata, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output [3:0]  io_out_bits_eccMask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
  output [3:0]  io_out_bits_way_en // @[:freechips.rocketchip.system.DefaultRV32Config.fir@115488.4]
);
  wire [3:0] _GEN_2; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115497.4]
  wire [31:0] _GEN_4; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115497.4]
  wire [11:0] _GEN_6; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115497.4]
  wire [3:0] _GEN_8; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  wire [3:0] _GEN_9; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  wire [31:0] _GEN_11; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  wire  _GEN_12; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  wire [11:0] _GEN_13; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  wire  _T; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@115524.4]
  wire  _T_1; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@115525.4]
  wire  _T_4; // @[Arbiter.scala 31:78:freechips.rocketchip.system.DefaultRV32Config.fir@115528.4]
  wire  _T_9; // @[Arbiter.scala 135:19:freechips.rocketchip.system.DefaultRV32Config.fir@115537.4]

  assign _GEN_2 = io_in_2_valid ? io_in_2_bits_eccMask : io_in_3_bits_eccMask; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115497.4]
  assign _GEN_4 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115497.4]
  assign _GEN_6 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115497.4]
  assign _GEN_8 = io_in_1_valid ? io_in_1_bits_way_en : 4'hf; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  assign _GEN_9 = io_in_1_valid ? 4'hf : _GEN_2; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  assign _GEN_11 = io_in_1_valid ? io_in_1_bits_wdata : _GEN_4; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  assign _GEN_12 = io_in_1_valid & io_in_1_bits_write; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  assign _GEN_13 = io_in_1_valid ? io_in_1_bits_addr : _GEN_6; // @[Arbiter.scala 126:27:freechips.rocketchip.system.DefaultRV32Config.fir@115506.4]
  assign _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@115524.4]
  assign _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@115525.4]
  assign _T_4 = _T_1 == 1'h0; // @[Arbiter.scala 31:78:freechips.rocketchip.system.DefaultRV32Config.fir@115528.4]
  assign _T_9 = _T_4 == 1'h0; // @[Arbiter.scala 135:19:freechips.rocketchip.system.DefaultRV32Config.fir@115537.4]
  assign io_in_1_ready = io_in_0_valid == 1'h0; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@115532.4]
  assign io_in_2_ready = _T == 1'h0; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@115534.4]
  assign io_in_3_ready = _T_1 == 1'h0; // @[Arbiter.scala 134:14:freechips.rocketchip.system.DefaultRV32Config.fir@115536.4]
  assign io_out_valid = _T_9 | io_in_3_valid; // @[Arbiter.scala 135:16:freechips.rocketchip.system.DefaultRV32Config.fir@115539.4]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_13; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@115496.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115504.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115513.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115522.6]
  assign io_out_bits_write = io_in_0_valid ? io_in_0_bits_write : _GEN_12; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@115495.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115503.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115512.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115521.6]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : _GEN_11; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@115494.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115502.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115511.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115520.6]
  assign io_out_bits_eccMask = io_in_0_valid ? io_in_0_bits_eccMask : _GEN_9; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@115492.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115500.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115509.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115518.6]
  assign io_out_bits_way_en = io_in_0_valid ? io_in_0_bits_way_en : _GEN_8; // @[Arbiter.scala 124:15:freechips.rocketchip.system.DefaultRV32Config.fir@115491.4 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115499.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115508.6 Arbiter.scala 128:19:freechips.rocketchip.system.DefaultRV32Config.fir@115517.6]
endmodule
`endif // ___3

