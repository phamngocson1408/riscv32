`include "include_module.v"
`ifdef __MemoryBus
module MemoryBus(
  input         clock,
  input         reset,
  input         auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_ready,
  output        auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_valid,
  output [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_id,
  output [31:0] auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_addr,
  output [7:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_len,
  output [2:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_size,
  output [1:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_burst,
  output        auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_lock,
  output [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_cache,
  output [2:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_prot,
  output [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_qos,
  input         auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_ready,
  output        auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_valid,
  output [31:0] auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_bits_data,
  output [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_bits_strb,
  output        auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_bits_last,
  output        auto_coupler_to_memory_controller_named_axi4_axi4yank_out_b_ready,
  input         auto_coupler_to_memory_controller_named_axi4_axi4yank_out_b_valid,
  input  [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_b_bits_id,
  input  [1:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_b_bits_resp,
  input         auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_ready,
  output        auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_valid,
  output [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_id,
  output [31:0] auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_addr,
  output [7:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_len,
  output [2:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_size,
  output [1:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_burst,
  output        auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_lock,
  output [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_cache,
  output [2:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_prot,
  output [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_qos,
  output        auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_ready,
  input         auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_valid,
  input  [3:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_bits_id,
  input  [31:0] auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_bits_data,
  input  [1:0]  auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_bits_resp,
  input         auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_bits_last,
  output        auto_coupler_from_coherence_manager_binder_in_a_ready,
  input         auto_coupler_from_coherence_manager_binder_in_a_valid,
  input  [2:0]  auto_coupler_from_coherence_manager_binder_in_a_bits_opcode,
  input  [2:0]  auto_coupler_from_coherence_manager_binder_in_a_bits_param,
  input  [2:0]  auto_coupler_from_coherence_manager_binder_in_a_bits_size,
  input  [1:0]  auto_coupler_from_coherence_manager_binder_in_a_bits_source,
  input  [31:0] auto_coupler_from_coherence_manager_binder_in_a_bits_address,
  input  [3:0]  auto_coupler_from_coherence_manager_binder_in_a_bits_mask,
  input  [31:0] auto_coupler_from_coherence_manager_binder_in_a_bits_data,
  input         auto_coupler_from_coherence_manager_binder_in_a_bits_corrupt,
  input         auto_coupler_from_coherence_manager_binder_in_d_ready,
  output        auto_coupler_from_coherence_manager_binder_in_d_valid,
  output [2:0]  auto_coupler_from_coherence_manager_binder_in_d_bits_opcode,
  output [2:0]  auto_coupler_from_coherence_manager_binder_in_d_bits_size,
  output [1:0]  auto_coupler_from_coherence_manager_binder_in_d_bits_source,
  output        auto_coupler_from_coherence_manager_binder_in_d_bits_denied,
  output [31:0] auto_coupler_from_coherence_manager_binder_in_d_bits_data,
  output        auto_coupler_from_coherence_manager_binder_in_d_bits_corrupt
);
  wire  memory_bus_xbar_clock;
  wire  memory_bus_xbar_reset;
  wire  memory_bus_xbar_auto_in_a_ready;
  wire  memory_bus_xbar_auto_in_a_valid;
  wire [2:0] memory_bus_xbar_auto_in_a_bits_opcode;
  wire [2:0] memory_bus_xbar_auto_in_a_bits_param;
  wire [2:0] memory_bus_xbar_auto_in_a_bits_size;
  wire [1:0] memory_bus_xbar_auto_in_a_bits_source;
  wire [31:0] memory_bus_xbar_auto_in_a_bits_address;
  wire [3:0] memory_bus_xbar_auto_in_a_bits_mask;
  wire [31:0] memory_bus_xbar_auto_in_a_bits_data;
  wire  memory_bus_xbar_auto_in_a_bits_corrupt;
  wire  memory_bus_xbar_auto_in_d_ready;
  wire  memory_bus_xbar_auto_in_d_valid;
  wire [2:0] memory_bus_xbar_auto_in_d_bits_opcode;
  wire [2:0] memory_bus_xbar_auto_in_d_bits_size;
  wire [1:0] memory_bus_xbar_auto_in_d_bits_source;
  wire  memory_bus_xbar_auto_in_d_bits_denied;
  wire [31:0] memory_bus_xbar_auto_in_d_bits_data;
  wire  memory_bus_xbar_auto_in_d_bits_corrupt;
  wire  memory_bus_xbar_auto_out_a_ready;
  wire  memory_bus_xbar_auto_out_a_valid;
  wire [2:0] memory_bus_xbar_auto_out_a_bits_opcode;
  wire [2:0] memory_bus_xbar_auto_out_a_bits_param;
  wire [2:0] memory_bus_xbar_auto_out_a_bits_size;
  wire [1:0] memory_bus_xbar_auto_out_a_bits_source;
  wire [31:0] memory_bus_xbar_auto_out_a_bits_address;
  wire [3:0] memory_bus_xbar_auto_out_a_bits_mask;
  wire [31:0] memory_bus_xbar_auto_out_a_bits_data;
  wire  memory_bus_xbar_auto_out_a_bits_corrupt;
  wire  memory_bus_xbar_auto_out_d_ready;
  wire  memory_bus_xbar_auto_out_d_valid;
  wire [2:0] memory_bus_xbar_auto_out_d_bits_opcode;
  wire [2:0] memory_bus_xbar_auto_out_d_bits_size;
  wire [1:0] memory_bus_xbar_auto_out_d_bits_source;
  wire  memory_bus_xbar_auto_out_d_bits_denied;
  wire [31:0] memory_bus_xbar_auto_out_d_bits_data;
  wire  memory_bus_xbar_auto_out_d_bits_corrupt;
  wire  coupler_from_coherence_manager_clock;
  wire  coupler_from_coherence_manager_reset;
  wire  coupler_from_coherence_manager_auto_binder_in_a_ready;
  wire  coupler_from_coherence_manager_auto_binder_in_a_valid;
  wire [2:0] coupler_from_coherence_manager_auto_binder_in_a_bits_opcode;
  wire [2:0] coupler_from_coherence_manager_auto_binder_in_a_bits_param;
  wire [2:0] coupler_from_coherence_manager_auto_binder_in_a_bits_size;
  wire [1:0] coupler_from_coherence_manager_auto_binder_in_a_bits_source;
  wire [31:0] coupler_from_coherence_manager_auto_binder_in_a_bits_address;
  wire [3:0] coupler_from_coherence_manager_auto_binder_in_a_bits_mask;
  wire [31:0] coupler_from_coherence_manager_auto_binder_in_a_bits_data;
  wire  coupler_from_coherence_manager_auto_binder_in_a_bits_corrupt;
  wire  coupler_from_coherence_manager_auto_binder_in_d_ready;
  wire  coupler_from_coherence_manager_auto_binder_in_d_valid;
  wire [2:0] coupler_from_coherence_manager_auto_binder_in_d_bits_opcode;
  wire [2:0] coupler_from_coherence_manager_auto_binder_in_d_bits_size;
  wire [1:0] coupler_from_coherence_manager_auto_binder_in_d_bits_source;
  wire  coupler_from_coherence_manager_auto_binder_in_d_bits_denied;
  wire [31:0] coupler_from_coherence_manager_auto_binder_in_d_bits_data;
  wire  coupler_from_coherence_manager_auto_binder_in_d_bits_corrupt;
  wire  coupler_from_coherence_manager_auto_binder_out_a_ready;
  wire  coupler_from_coherence_manager_auto_binder_out_a_valid;
  wire [2:0] coupler_from_coherence_manager_auto_binder_out_a_bits_opcode;
  wire [2:0] coupler_from_coherence_manager_auto_binder_out_a_bits_param;
  wire [2:0] coupler_from_coherence_manager_auto_binder_out_a_bits_size;
  wire [1:0] coupler_from_coherence_manager_auto_binder_out_a_bits_source;
  wire [31:0] coupler_from_coherence_manager_auto_binder_out_a_bits_address;
  wire [3:0] coupler_from_coherence_manager_auto_binder_out_a_bits_mask;
  wire [31:0] coupler_from_coherence_manager_auto_binder_out_a_bits_data;
  wire  coupler_from_coherence_manager_auto_binder_out_a_bits_corrupt;
  wire  coupler_from_coherence_manager_auto_binder_out_d_ready;
  wire  coupler_from_coherence_manager_auto_binder_out_d_valid;
  wire [2:0] coupler_from_coherence_manager_auto_binder_out_d_bits_opcode;
  wire [2:0] coupler_from_coherence_manager_auto_binder_out_d_bits_size;
  wire [1:0] coupler_from_coherence_manager_auto_binder_out_d_bits_source;
  wire  coupler_from_coherence_manager_auto_binder_out_d_bits_denied;
  wire [31:0] coupler_from_coherence_manager_auto_binder_out_d_bits_data;
  wire  coupler_from_coherence_manager_auto_binder_out_d_bits_corrupt;
  wire  coupler_to_memory_controller_named_axi4_clock;
  wire  coupler_to_memory_controller_named_axi4_reset;
  wire  coupler_to_memory_controller_named_axi4_auto_picker_in_a_ready;
  wire  coupler_to_memory_controller_named_axi4_auto_picker_in_a_valid;
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_opcode;
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_param;
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_size;
  wire [1:0] coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_source;
  wire [31:0] coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_address;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_mask;
  wire [31:0] coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_data;
  wire  coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_corrupt;
  wire  coupler_to_memory_controller_named_axi4_auto_picker_in_d_ready;
  wire  coupler_to_memory_controller_named_axi4_auto_picker_in_d_valid;
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_opcode;
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_size;
  wire [1:0] coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_source;
  wire  coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_denied;
  wire [31:0] coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_data;
  wire  coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_corrupt;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_ready;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_valid;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_id;
  wire [31:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_addr;
  wire [7:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_len;
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_size;
  wire [1:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_burst;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_lock;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_cache;
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_prot;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_qos;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_ready;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_valid;
  wire [31:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_data;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_strb;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_last; 
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_ready;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_valid;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_bits_id;
  wire [1:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_bits_resp;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_ready;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_valid;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_id;
  wire [31:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_addr;
  wire [7:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_len; 
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_size; 
  wire [1:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_burst;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_lock;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_cache; 
  wire [2:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_prot;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_qos;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_ready;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_valid;
  wire [3:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_id;
  wire [31:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_data; 
  wire [1:0] coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_resp;
  wire  coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_last; 
  TLXbar_4 memory_bus_xbar (
    .clock(memory_bus_xbar_clock),
    .reset(memory_bus_xbar_reset),
    .auto_in_a_ready(memory_bus_xbar_auto_in_a_ready),
    .auto_in_a_valid(memory_bus_xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(memory_bus_xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(memory_bus_xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(memory_bus_xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(memory_bus_xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(memory_bus_xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(memory_bus_xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(memory_bus_xbar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(memory_bus_xbar_auto_in_a_bits_corrupt),
    .auto_in_d_ready(memory_bus_xbar_auto_in_d_ready),
    .auto_in_d_valid(memory_bus_xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(memory_bus_xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(memory_bus_xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(memory_bus_xbar_auto_in_d_bits_source),
    .auto_in_d_bits_denied(memory_bus_xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(memory_bus_xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(memory_bus_xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(memory_bus_xbar_auto_out_a_ready),
    .auto_out_a_valid(memory_bus_xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(memory_bus_xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(memory_bus_xbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(memory_bus_xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(memory_bus_xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(memory_bus_xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(memory_bus_xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(memory_bus_xbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(memory_bus_xbar_auto_out_a_bits_corrupt),
    .auto_out_d_ready(memory_bus_xbar_auto_out_d_ready),
    .auto_out_d_valid(memory_bus_xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(memory_bus_xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(memory_bus_xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(memory_bus_xbar_auto_out_d_bits_source),
    .auto_out_d_bits_denied(memory_bus_xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(memory_bus_xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(memory_bus_xbar_auto_out_d_bits_corrupt)
  );
  SimpleLazyModule_6 coupler_from_coherence_manager ( 
    .clock(coupler_from_coherence_manager_clock),
    .reset(coupler_from_coherence_manager_reset),
    .auto_binder_in_a_ready(coupler_from_coherence_manager_auto_binder_in_a_ready),
    .auto_binder_in_a_valid(coupler_from_coherence_manager_auto_binder_in_a_valid),
    .auto_binder_in_a_bits_opcode(coupler_from_coherence_manager_auto_binder_in_a_bits_opcode),
    .auto_binder_in_a_bits_param(coupler_from_coherence_manager_auto_binder_in_a_bits_param),
    .auto_binder_in_a_bits_size(coupler_from_coherence_manager_auto_binder_in_a_bits_size),
    .auto_binder_in_a_bits_source(coupler_from_coherence_manager_auto_binder_in_a_bits_source),
    .auto_binder_in_a_bits_address(coupler_from_coherence_manager_auto_binder_in_a_bits_address),
    .auto_binder_in_a_bits_mask(coupler_from_coherence_manager_auto_binder_in_a_bits_mask),
    .auto_binder_in_a_bits_data(coupler_from_coherence_manager_auto_binder_in_a_bits_data),
    .auto_binder_in_a_bits_corrupt(coupler_from_coherence_manager_auto_binder_in_a_bits_corrupt),
    .auto_binder_in_d_ready(coupler_from_coherence_manager_auto_binder_in_d_ready),
    .auto_binder_in_d_valid(coupler_from_coherence_manager_auto_binder_in_d_valid),
    .auto_binder_in_d_bits_opcode(coupler_from_coherence_manager_auto_binder_in_d_bits_opcode),
    .auto_binder_in_d_bits_size(coupler_from_coherence_manager_auto_binder_in_d_bits_size),
    .auto_binder_in_d_bits_source(coupler_from_coherence_manager_auto_binder_in_d_bits_source),
    .auto_binder_in_d_bits_denied(coupler_from_coherence_manager_auto_binder_in_d_bits_denied),
    .auto_binder_in_d_bits_data(coupler_from_coherence_manager_auto_binder_in_d_bits_data),
    .auto_binder_in_d_bits_corrupt(coupler_from_coherence_manager_auto_binder_in_d_bits_corrupt),
    .auto_binder_out_a_ready(coupler_from_coherence_manager_auto_binder_out_a_ready),
    .auto_binder_out_a_valid(coupler_from_coherence_manager_auto_binder_out_a_valid),
    .auto_binder_out_a_bits_opcode(coupler_from_coherence_manager_auto_binder_out_a_bits_opcode),
    .auto_binder_out_a_bits_param(coupler_from_coherence_manager_auto_binder_out_a_bits_param),
    .auto_binder_out_a_bits_size(coupler_from_coherence_manager_auto_binder_out_a_bits_size),
    .auto_binder_out_a_bits_source(coupler_from_coherence_manager_auto_binder_out_a_bits_source),
    .auto_binder_out_a_bits_address(coupler_from_coherence_manager_auto_binder_out_a_bits_address),
    .auto_binder_out_a_bits_mask(coupler_from_coherence_manager_auto_binder_out_a_bits_mask),
    .auto_binder_out_a_bits_data(coupler_from_coherence_manager_auto_binder_out_a_bits_data),
    .auto_binder_out_a_bits_corrupt(coupler_from_coherence_manager_auto_binder_out_a_bits_corrupt),
    .auto_binder_out_d_ready(coupler_from_coherence_manager_auto_binder_out_d_ready),
    .auto_binder_out_d_valid(coupler_from_coherence_manager_auto_binder_out_d_valid),
    .auto_binder_out_d_bits_opcode(coupler_from_coherence_manager_auto_binder_out_d_bits_opcode),
    .auto_binder_out_d_bits_size(coupler_from_coherence_manager_auto_binder_out_d_bits_size),
    .auto_binder_out_d_bits_source(coupler_from_coherence_manager_auto_binder_out_d_bits_source),
    .auto_binder_out_d_bits_denied(coupler_from_coherence_manager_auto_binder_out_d_bits_denied),
    .auto_binder_out_d_bits_data(coupler_from_coherence_manager_auto_binder_out_d_bits_data),
    .auto_binder_out_d_bits_corrupt(coupler_from_coherence_manager_auto_binder_out_d_bits_corrupt)
  );
  SimpleLazyModule_7 coupler_to_memory_controller_named_axi4 (
    .clock(coupler_to_memory_controller_named_axi4_clock),
    .reset(coupler_to_memory_controller_named_axi4_reset),
    .auto_picker_in_a_ready(coupler_to_memory_controller_named_axi4_auto_picker_in_a_ready),
    .auto_picker_in_a_valid(coupler_to_memory_controller_named_axi4_auto_picker_in_a_valid),
    .auto_picker_in_a_bits_opcode(coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_opcode),
    .auto_picker_in_a_bits_param(coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_param),
    .auto_picker_in_a_bits_size(coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_size),
    .auto_picker_in_a_bits_source(coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_source),
    .auto_picker_in_a_bits_address(coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_address),
    .auto_picker_in_a_bits_mask(coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_mask),
    .auto_picker_in_a_bits_data(coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_data),
    .auto_picker_in_a_bits_corrupt(coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_corrupt),
    .auto_picker_in_d_ready(coupler_to_memory_controller_named_axi4_auto_picker_in_d_ready),
    .auto_picker_in_d_valid(coupler_to_memory_controller_named_axi4_auto_picker_in_d_valid),
    .auto_picker_in_d_bits_opcode(coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_opcode),
    .auto_picker_in_d_bits_size(coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_size),
    .auto_picker_in_d_bits_source(coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_source),
    .auto_picker_in_d_bits_denied(coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_denied),
    .auto_picker_in_d_bits_data(coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_data),
    .auto_picker_in_d_bits_corrupt(coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_corrupt),
    .auto_axi4yank_out_aw_ready(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_ready),
    .auto_axi4yank_out_aw_valid(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_valid),
    .auto_axi4yank_out_aw_bits_id(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_id),
    .auto_axi4yank_out_aw_bits_addr(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_addr),
    .auto_axi4yank_out_aw_bits_len(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_len),
    .auto_axi4yank_out_aw_bits_size(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_size),
    .auto_axi4yank_out_aw_bits_burst(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_burst),
    .auto_axi4yank_out_aw_bits_lock(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_lock),
    .auto_axi4yank_out_aw_bits_cache(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_cache),
    .auto_axi4yank_out_aw_bits_prot(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_prot),
    .auto_axi4yank_out_aw_bits_qos(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_qos),
    .auto_axi4yank_out_w_ready(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_ready),
    .auto_axi4yank_out_w_valid(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_valid),
    .auto_axi4yank_out_w_bits_data(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_data),
    .auto_axi4yank_out_w_bits_strb(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_strb),
    .auto_axi4yank_out_w_bits_last(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_last),
    .auto_axi4yank_out_b_ready(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_ready),
    .auto_axi4yank_out_b_valid(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_valid),
    .auto_axi4yank_out_b_bits_id(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_bits_id),
    .auto_axi4yank_out_b_bits_resp(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_bits_resp),
    .auto_axi4yank_out_ar_ready(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_ready),
    .auto_axi4yank_out_ar_valid(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_valid),
    .auto_axi4yank_out_ar_bits_id(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_id),
    .auto_axi4yank_out_ar_bits_addr(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_addr),
    .auto_axi4yank_out_ar_bits_len(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_len),
    .auto_axi4yank_out_ar_bits_size(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_size),
    .auto_axi4yank_out_ar_bits_burst(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_burst),
    .auto_axi4yank_out_ar_bits_lock(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_lock),
    .auto_axi4yank_out_ar_bits_cache(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_cache),
    .auto_axi4yank_out_ar_bits_prot(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_prot),
    .auto_axi4yank_out_ar_bits_qos(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_qos),
    .auto_axi4yank_out_r_ready(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_ready),
    .auto_axi4yank_out_r_valid(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_valid),
    .auto_axi4yank_out_r_bits_id(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_id),
    .auto_axi4yank_out_r_bits_data(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_data),
    .auto_axi4yank_out_r_bits_resp(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_resp),
    .auto_axi4yank_out_r_bits_last(coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_last)
  );
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_valid = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_valid;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_id = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_id;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_addr = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_addr;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_len = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_len; 
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_size = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_size;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_burst = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_burst;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_lock = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_lock;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_cache = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_cache;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_prot = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_prot;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_bits_qos = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_bits_qos;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_valid = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_valid;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_bits_data = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_data;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_bits_strb = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_strb;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_bits_last = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_bits_last;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_b_ready = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_ready; 
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_valid = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_valid;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_id = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_id;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_addr = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_addr;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_len = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_len;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_size = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_size;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_burst = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_burst;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_lock = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_lock;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_cache = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_cache;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_prot = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_prot;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_bits_qos = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_bits_qos;
  assign auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_ready = coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_ready; 
  assign auto_coupler_from_coherence_manager_binder_in_a_ready = coupler_from_coherence_manager_auto_binder_in_a_ready;
  assign auto_coupler_from_coherence_manager_binder_in_d_valid = coupler_from_coherence_manager_auto_binder_in_d_valid;
  assign auto_coupler_from_coherence_manager_binder_in_d_bits_opcode = coupler_from_coherence_manager_auto_binder_in_d_bits_opcode;
  assign auto_coupler_from_coherence_manager_binder_in_d_bits_size = coupler_from_coherence_manager_auto_binder_in_d_bits_size; 
  assign auto_coupler_from_coherence_manager_binder_in_d_bits_source = coupler_from_coherence_manager_auto_binder_in_d_bits_source; 
  assign auto_coupler_from_coherence_manager_binder_in_d_bits_denied = coupler_from_coherence_manager_auto_binder_in_d_bits_denied;
  assign auto_coupler_from_coherence_manager_binder_in_d_bits_data = coupler_from_coherence_manager_auto_binder_in_d_bits_data;
  assign auto_coupler_from_coherence_manager_binder_in_d_bits_corrupt = coupler_from_coherence_manager_auto_binder_in_d_bits_corrupt;
  assign memory_bus_xbar_clock = clock;
  assign memory_bus_xbar_reset = reset;
  assign memory_bus_xbar_auto_in_a_valid = coupler_from_coherence_manager_auto_binder_out_a_valid;
  assign memory_bus_xbar_auto_in_a_bits_opcode = coupler_from_coherence_manager_auto_binder_out_a_bits_opcode;
  assign memory_bus_xbar_auto_in_a_bits_param = coupler_from_coherence_manager_auto_binder_out_a_bits_param;
  assign memory_bus_xbar_auto_in_a_bits_size = coupler_from_coherence_manager_auto_binder_out_a_bits_size; 
  assign memory_bus_xbar_auto_in_a_bits_source = coupler_from_coherence_manager_auto_binder_out_a_bits_source;
  assign memory_bus_xbar_auto_in_a_bits_address = coupler_from_coherence_manager_auto_binder_out_a_bits_address;
  assign memory_bus_xbar_auto_in_a_bits_mask = coupler_from_coherence_manager_auto_binder_out_a_bits_mask; 
  assign memory_bus_xbar_auto_in_a_bits_data = coupler_from_coherence_manager_auto_binder_out_a_bits_data; 
  assign memory_bus_xbar_auto_in_a_bits_corrupt = coupler_from_coherence_manager_auto_binder_out_a_bits_corrupt;
  assign memory_bus_xbar_auto_in_d_ready = coupler_from_coherence_manager_auto_binder_out_d_ready;
  assign memory_bus_xbar_auto_out_a_ready = coupler_to_memory_controller_named_axi4_auto_picker_in_a_ready; 
  assign memory_bus_xbar_auto_out_d_valid = coupler_to_memory_controller_named_axi4_auto_picker_in_d_valid;
  assign memory_bus_xbar_auto_out_d_bits_opcode = coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_opcode;
  assign memory_bus_xbar_auto_out_d_bits_size = coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_size;
  assign memory_bus_xbar_auto_out_d_bits_source = coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_source;
  assign memory_bus_xbar_auto_out_d_bits_denied = coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_denied;
  assign memory_bus_xbar_auto_out_d_bits_data = coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_data;
  assign memory_bus_xbar_auto_out_d_bits_corrupt = coupler_to_memory_controller_named_axi4_auto_picker_in_d_bits_corrupt;
  assign coupler_from_coherence_manager_clock = clock;
  assign coupler_from_coherence_manager_reset = reset;
  assign coupler_from_coherence_manager_auto_binder_in_a_valid = auto_coupler_from_coherence_manager_binder_in_a_valid;
  assign coupler_from_coherence_manager_auto_binder_in_a_bits_opcode = auto_coupler_from_coherence_manager_binder_in_a_bits_opcode;
  assign coupler_from_coherence_manager_auto_binder_in_a_bits_param = auto_coupler_from_coherence_manager_binder_in_a_bits_param;
  assign coupler_from_coherence_manager_auto_binder_in_a_bits_size = auto_coupler_from_coherence_manager_binder_in_a_bits_size; 
  assign coupler_from_coherence_manager_auto_binder_in_a_bits_source = auto_coupler_from_coherence_manager_binder_in_a_bits_source;
  assign coupler_from_coherence_manager_auto_binder_in_a_bits_address = auto_coupler_from_coherence_manager_binder_in_a_bits_address;
  assign coupler_from_coherence_manager_auto_binder_in_a_bits_mask = auto_coupler_from_coherence_manager_binder_in_a_bits_mask;
  assign coupler_from_coherence_manager_auto_binder_in_a_bits_data = auto_coupler_from_coherence_manager_binder_in_a_bits_data;
  assign coupler_from_coherence_manager_auto_binder_in_a_bits_corrupt = auto_coupler_from_coherence_manager_binder_in_a_bits_corrupt;
  assign coupler_from_coherence_manager_auto_binder_in_d_ready = auto_coupler_from_coherence_manager_binder_in_d_ready;
  assign coupler_from_coherence_manager_auto_binder_out_a_ready = memory_bus_xbar_auto_in_a_ready;
  assign coupler_from_coherence_manager_auto_binder_out_d_valid = memory_bus_xbar_auto_in_d_valid; 
  assign coupler_from_coherence_manager_auto_binder_out_d_bits_opcode = memory_bus_xbar_auto_in_d_bits_opcode;
  assign coupler_from_coherence_manager_auto_binder_out_d_bits_size = memory_bus_xbar_auto_in_d_bits_size;
  assign coupler_from_coherence_manager_auto_binder_out_d_bits_source = memory_bus_xbar_auto_in_d_bits_source;
  assign coupler_from_coherence_manager_auto_binder_out_d_bits_denied = memory_bus_xbar_auto_in_d_bits_denied;
  assign coupler_from_coherence_manager_auto_binder_out_d_bits_data = memory_bus_xbar_auto_in_d_bits_data;
  assign coupler_from_coherence_manager_auto_binder_out_d_bits_corrupt = memory_bus_xbar_auto_in_d_bits_corrupt;
  assign coupler_to_memory_controller_named_axi4_clock = clock;
  assign coupler_to_memory_controller_named_axi4_reset = reset;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_valid = memory_bus_xbar_auto_out_a_valid;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_opcode = memory_bus_xbar_auto_out_a_bits_opcode;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_param = memory_bus_xbar_auto_out_a_bits_param;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_size = memory_bus_xbar_auto_out_a_bits_size;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_source = memory_bus_xbar_auto_out_a_bits_source;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_address = memory_bus_xbar_auto_out_a_bits_address;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_mask = memory_bus_xbar_auto_out_a_bits_mask;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_data = memory_bus_xbar_auto_out_a_bits_data;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_a_bits_corrupt = memory_bus_xbar_auto_out_a_bits_corrupt;
  assign coupler_to_memory_controller_named_axi4_auto_picker_in_d_ready = memory_bus_xbar_auto_out_d_ready;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_aw_ready = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_aw_ready;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_w_ready = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_w_ready;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_valid = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_b_valid;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_bits_id = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_b_bits_id;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_b_bits_resp = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_b_bits_resp;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_ar_ready = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_ar_ready;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_valid = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_valid;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_id = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_bits_id;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_data = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_bits_data;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_resp = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_bits_resp;
  assign coupler_to_memory_controller_named_axi4_auto_axi4yank_out_r_bits_last = auto_coupler_to_memory_controller_named_axi4_axi4yank_out_r_bits_last;
endmodule
`endif // __MemoryBus

