`include "include_module.v"
`ifdef __CSRFile
module CSRFile( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170045.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170046.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170047.4]
  input         io_ungated_clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input         io_interrupts_debug, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input         io_interrupts_mtip, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input         io_interrupts_msip, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input         io_interrupts_meip, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [11:0] io_rw_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [2:0]  io_rw_cmd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_rw_rdata, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [31:0] io_rw_wdata, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [11:0] io_decode_0_csr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_decode_0_fp_illegal, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_decode_0_fp_csr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_decode_0_read_illegal, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_decode_0_write_illegal, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_decode_0_write_flush, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_decode_0_system_illegal, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_csr_stall, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_eret, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_singleStep, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_debug, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_cease, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_status_isa, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_dprv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_prv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_sd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [26:0] io_status_zero2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_sxl, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_uxl, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_sd_rv32, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [5:0]  io_status_zero1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_vs, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_tsr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_tw, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_tvm, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_mxr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_sum, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_mprv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_xs, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_fs, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_mpp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_status_hpp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_spp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_mpie, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_hpie, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_spie, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_upie, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_mie, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_hie, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_sie, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_status_uie, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_evec, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input         io_exception, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input         io_retire, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [31:0] io_cause, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [31:0] io_pc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [31:0] io_tval, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_time, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [2:0]  io_fcsr_rm, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input         io_fcsr_flags_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [4:0]  io_fcsr_flags_bits, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_interrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_interrupt_cause, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_bp_0_control_action, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_bp_0_control_tmatch, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_bp_0_control_m, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_bp_0_control_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_bp_0_control_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_bp_0_control_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_bp_0_control_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_bp_0_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_0_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_pmp_0_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_0_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_0_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_0_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [29:0] io_pmp_0_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_pmp_0_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_1_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_pmp_1_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_1_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_1_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_1_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [29:0] io_pmp_1_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_pmp_1_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_2_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_pmp_2_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_2_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_2_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_2_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [29:0] io_pmp_2_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_pmp_2_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_3_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_pmp_3_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_3_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_3_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_3_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [29:0] io_pmp_3_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_pmp_3_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_4_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_pmp_4_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_4_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_4_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_4_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [29:0] io_pmp_4_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_pmp_4_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_5_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_pmp_5_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_5_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_5_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_5_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [29:0] io_pmp_5_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_pmp_5_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_6_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_pmp_6_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_6_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_6_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_6_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [29:0] io_pmp_6_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_pmp_6_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_7_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [1:0]  io_pmp_7_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_7_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_7_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_pmp_7_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [29:0] io_pmp_7_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_pmp_7_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  input  [31:0] io_inst_0, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_trace_0_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_trace_0_iaddr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output [31:0] io_trace_0_insn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
  output        io_trace_0_exception // @[:freechips.rocketchip.system.DefaultRV32Config.fir@170048.4]
);
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 299:24:freechips.rocketchip.system.DefaultRV32Config.fir@170125.4]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_mprv; // @[CSR.scala 299:24:freechips.rocketchip.system.DefaultRV32Config.fir@170125.4]
  reg [31:0] _RAND_1;
  reg [1:0] reg_mstatus_fs; // @[CSR.scala 299:24:freechips.rocketchip.system.DefaultRV32Config.fir@170125.4]
  reg [31:0] _RAND_2;
  reg [1:0] reg_mstatus_mpp; // @[CSR.scala 299:24:freechips.rocketchip.system.DefaultRV32Config.fir@170125.4]
  reg [31:0] _RAND_3;
  reg  reg_mstatus_spp; // @[CSR.scala 299:24:freechips.rocketchip.system.DefaultRV32Config.fir@170125.4]
  reg [31:0] _RAND_4;
  reg  reg_mstatus_mpie; // @[CSR.scala 299:24:freechips.rocketchip.system.DefaultRV32Config.fir@170125.4]
  reg [31:0] _RAND_5;
  reg  reg_mstatus_mie; // @[CSR.scala 299:24:freechips.rocketchip.system.DefaultRV32Config.fir@170125.4]
  reg [31:0] _RAND_6;
  wire  system_insn; // @[CSR.scala 574:31:freechips.rocketchip.system.DefaultRV32Config.fir@171058.4]
  wire [31:0] _T_804; // @[CSR.scala 586:28:freechips.rocketchip.system.DefaultRV32Config.fir@171059.4]
  wire [31:0] _T_811; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171066.4]
  wire  _T_812; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171067.4]
  wire  insn_ret; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171080.4]
  wire  _T_1729; // @[CSR.scala 729:47:freechips.rocketchip.system.DefaultRV32Config.fir@172091.8]
  reg [1:0] reg_dcsr_prv; // @[CSR.scala 307:21:freechips.rocketchip.system.DefaultRV32Config.fir@170171.4]
  reg [31:0] _RAND_7;
  wire [1:0] _GEN_93; // @[CSR.scala 729:53:freechips.rocketchip.system.DefaultRV32Config.fir@172093.8]
  wire [31:0] _T_805; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171060.4]
  wire  _T_806; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171061.4]
  wire  insn_call; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171076.4]
  wire [31:0] _T_808; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171063.4]
  wire  _T_809; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171064.4]
  wire  insn_break; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171078.4]
  wire  _T_1388; // @[CSR.scala 658:29:freechips.rocketchip.system.DefaultRV32Config.fir@171680.4]
  wire  exception; // @[CSR.scala 658:43:freechips.rocketchip.system.DefaultRV32Config.fir@171681.4]
  reg  reg_singleStepped; // @[CSR.scala 351:30:freechips.rocketchip.system.DefaultRV32Config.fir@170230.4]
  reg [31:0] _RAND_8;
  wire [3:0] _GEN_439; // @[CSR.scala 622:36:freechips.rocketchip.system.DefaultRV32Config.fir@171602.4]
  wire [3:0] _T_1334; // @[CSR.scala 622:36:freechips.rocketchip.system.DefaultRV32Config.fir@171603.4]
  wire [31:0] _T_1335; // @[CSR.scala 623:14:freechips.rocketchip.system.DefaultRV32Config.fir@171604.4]
  wire [31:0] cause; // @[CSR.scala 622:8:freechips.rocketchip.system.DefaultRV32Config.fir@171605.4]
  wire  _T_1336; // @[CSR.scala 625:30:freechips.rocketchip.system.DefaultRV32Config.fir@171607.4]
  wire [7:0] cause_lsbs; // @[CSR.scala 624:25:freechips.rocketchip.system.DefaultRV32Config.fir@171606.4]
  wire  _T_1337; // @[CSR.scala 625:53:freechips.rocketchip.system.DefaultRV32Config.fir@171608.4]
  wire  causeIsDebugInt; // @[CSR.scala 625:39:freechips.rocketchip.system.DefaultRV32Config.fir@171609.4]
  wire  _T_1349; // @[CSR.scala 628:60:freechips.rocketchip.system.DefaultRV32Config.fir@171623.4]
  wire  _T_1339; // @[CSR.scala 626:29:freechips.rocketchip.system.DefaultRV32Config.fir@171611.4]
  wire  causeIsDebugTrigger; // @[CSR.scala 626:44:freechips.rocketchip.system.DefaultRV32Config.fir@171613.4]
  wire  _T_1350; // @[CSR.scala 628:79:freechips.rocketchip.system.DefaultRV32Config.fir@171624.4]
  wire  _T_1343; // @[CSR.scala 627:42:freechips.rocketchip.system.DefaultRV32Config.fir@171616.4]
  reg  reg_dcsr_ebreakm; // @[CSR.scala 307:21:freechips.rocketchip.system.DefaultRV32Config.fir@170171.4]
  reg [31:0] _RAND_9;
  reg  reg_dcsr_ebreaku; // @[CSR.scala 307:21:freechips.rocketchip.system.DefaultRV32Config.fir@170171.4]
  reg [31:0] _RAND_10;
  wire [3:0] _T_1346; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@171619.4]
  wire [3:0] _T_1347; // @[CSR.scala 627:134:freechips.rocketchip.system.DefaultRV32Config.fir@171620.4]
  wire  _T_1348; // @[CSR.scala 627:134:freechips.rocketchip.system.DefaultRV32Config.fir@171621.4]
  wire  causeIsDebugBreak; // @[CSR.scala 627:56:freechips.rocketchip.system.DefaultRV32Config.fir@171622.4]
  wire  _T_1351; // @[CSR.scala 628:102:freechips.rocketchip.system.DefaultRV32Config.fir@171625.4]
  reg  reg_debug; // @[CSR.scala 348:22:freechips.rocketchip.system.DefaultRV32Config.fir@170227.4]
  reg [31:0] _RAND_11;
  wire  trapToDebug; // @[CSR.scala 628:123:freechips.rocketchip.system.DefaultRV32Config.fir@171626.4]
  wire  _T_1423; // @[CSR.scala 675:13:freechips.rocketchip.system.DefaultRV32Config.fir@171746.8]
  wire [1:0] _GEN_42; // @[CSR.scala 675:25:freechips.rocketchip.system.DefaultRV32Config.fir@171747.8]
  wire  _T_1354; // @[CSR.scala 630:51:freechips.rocketchip.system.DefaultRV32Config.fir@171630.4]
  wire [1:0] _GEN_61; // @[CSR.scala 674:24:freechips.rocketchip.system.DefaultRV32Config.fir@171745.6]
  wire [1:0] _GEN_79; // @[CSR.scala 673:20:freechips.rocketchip.system.DefaultRV32Config.fir@171744.4]
  wire [1:0] new_prv; // @[CSR.scala 722:19:freechips.rocketchip.system.DefaultRV32Config.fir@172074.4]
  wire  _T_33; // @[CSR.scala 1048:37:freechips.rocketchip.system.DefaultRV32Config.fir@170129.4]
  reg [2:0] reg_dcsr_cause; // @[CSR.scala 307:21:freechips.rocketchip.system.DefaultRV32Config.fir@170171.4]
  reg [31:0] _RAND_12;
  reg  reg_dcsr_step; // @[CSR.scala 307:21:freechips.rocketchip.system.DefaultRV32Config.fir@170171.4]
  reg [31:0] _RAND_13;
  reg [31:0] reg_dpc; // @[CSR.scala 349:20:freechips.rocketchip.system.DefaultRV32Config.fir@170228.4]
  reg [31:0] _RAND_14;
  reg [31:0] reg_dscratch; // @[CSR.scala 350:25:freechips.rocketchip.system.DefaultRV32Config.fir@170229.4]
  reg [31:0] _RAND_15;
  reg  reg_bp_0_control_dmode; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_16;
  reg  reg_bp_0_control_action; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_17;
  reg [1:0] reg_bp_0_control_tmatch; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_18;
  reg  reg_bp_0_control_m; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_19;
  reg  reg_bp_0_control_u; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_20;
  reg  reg_bp_0_control_x; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_21;
  reg  reg_bp_0_control_w; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_22;
  reg  reg_bp_0_control_r; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_23;
  reg [31:0] reg_bp_0_address; // @[CSR.scala 354:19:freechips.rocketchip.system.DefaultRV32Config.fir@170232.4]
  reg [31:0] _RAND_24;
  reg  reg_pmp_0_cfg_l; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_25;
  reg [1:0] reg_pmp_0_cfg_a; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_26;
  reg  reg_pmp_0_cfg_x; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_27;
  reg  reg_pmp_0_cfg_w; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_28;
  reg  reg_pmp_0_cfg_r; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_29;
  reg [29:0] reg_pmp_0_addr; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_30;
  reg  reg_pmp_1_cfg_l; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_31;
  reg [1:0] reg_pmp_1_cfg_a; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_32;
  reg  reg_pmp_1_cfg_x; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_33;
  reg  reg_pmp_1_cfg_w; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_34;
  reg  reg_pmp_1_cfg_r; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_35;
  reg [29:0] reg_pmp_1_addr; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_36;
  reg  reg_pmp_2_cfg_l; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_37;
  reg [1:0] reg_pmp_2_cfg_a; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_38;
  reg  reg_pmp_2_cfg_x; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_39;
  reg  reg_pmp_2_cfg_w; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_40;
  reg  reg_pmp_2_cfg_r; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_41;
  reg [29:0] reg_pmp_2_addr; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_42;
  reg  reg_pmp_3_cfg_l; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_43;
  reg [1:0] reg_pmp_3_cfg_a; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_44;
  reg  reg_pmp_3_cfg_x; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_45;
  reg  reg_pmp_3_cfg_w; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_46;
  reg  reg_pmp_3_cfg_r; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_47;
  reg [29:0] reg_pmp_3_addr; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_48;
  reg  reg_pmp_4_cfg_l; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_49;
  reg [1:0] reg_pmp_4_cfg_a; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_50;
  reg  reg_pmp_4_cfg_x; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_51;
  reg  reg_pmp_4_cfg_w; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_52;
  reg  reg_pmp_4_cfg_r; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_53;
  reg [29:0] reg_pmp_4_addr; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_54;
  reg  reg_pmp_5_cfg_l; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_55;
  reg [1:0] reg_pmp_5_cfg_a; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_56;
  reg  reg_pmp_5_cfg_x; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_57;
  reg  reg_pmp_5_cfg_w; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_58;
  reg  reg_pmp_5_cfg_r; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_59;
  reg [29:0] reg_pmp_5_addr; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_60;
  reg  reg_pmp_6_cfg_l; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_61;
  reg [1:0] reg_pmp_6_cfg_a; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_62;
  reg  reg_pmp_6_cfg_x; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_63;
  reg  reg_pmp_6_cfg_w; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_64;
  reg  reg_pmp_6_cfg_r; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_65;
  reg [29:0] reg_pmp_6_addr; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_66;
  reg  reg_pmp_7_cfg_l; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_67;
  reg [1:0] reg_pmp_7_cfg_a; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_68;
  reg  reg_pmp_7_cfg_x; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_69;
  reg  reg_pmp_7_cfg_w; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_70;
  reg  reg_pmp_7_cfg_r; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_71;
  reg [29:0] reg_pmp_7_addr; // @[CSR.scala 355:20:freechips.rocketchip.system.DefaultRV32Config.fir@170233.4]
  reg [31:0] _RAND_72;
  reg [31:0] reg_mie; // @[CSR.scala 357:20:freechips.rocketchip.system.DefaultRV32Config.fir@170234.4]
  reg [31:0] _RAND_73;
  reg [31:0] reg_mepc; // @[CSR.scala 367:21:freechips.rocketchip.system.DefaultRV32Config.fir@170242.4]
  reg [31:0] _RAND_74;
  reg [31:0] reg_mcause; // @[CSR.scala 368:23:freechips.rocketchip.system.DefaultRV32Config.fir@170243.4]
  reg [31:0] _RAND_75;
  reg [31:0] reg_mtval; // @[CSR.scala 369:22:freechips.rocketchip.system.DefaultRV32Config.fir@170244.4]
  reg [31:0] _RAND_76;
  reg [31:0] reg_mscratch; // @[CSR.scala 370:25:freechips.rocketchip.system.DefaultRV32Config.fir@170245.4]
  reg [31:0] _RAND_77;
  reg [31:0] reg_mtvec; // @[CSR.scala 373:27:freechips.rocketchip.system.DefaultRV32Config.fir@170246.4]
  reg [31:0] _RAND_78;
  reg [31:0] reg_mcounteren; // @[CSR.scala 379:18:freechips.rocketchip.system.DefaultRV32Config.fir@170247.4]
  reg [31:0] _RAND_79;
  wire [31:0] read_mcounteren; // @[CSR.scala 380:30:freechips.rocketchip.system.DefaultRV32Config.fir@170248.4]
  reg  reg_wfi; // @[CSR.scala 393:50:freechips.rocketchip.system.DefaultRV32Config.fir@170259.4]
  reg [31:0] _RAND_80;
  reg [4:0] reg_fflags; // @[CSR.scala 395:23:freechips.rocketchip.system.DefaultRV32Config.fir@170260.4]
  reg [31:0] _RAND_81;
  reg [2:0] reg_frm; // @[CSR.scala 396:20:freechips.rocketchip.system.DefaultRV32Config.fir@170261.4]
  reg [31:0] _RAND_82;
  reg [5:0] _T_87; // @[Counters.scala 46:37:freechips.rocketchip.system.DefaultRV32Config.fir@170262.4]
  reg [31:0] _RAND_83;
  wire [5:0] _GEN_440; // @[Counters.scala 47:33:freechips.rocketchip.system.DefaultRV32Config.fir@170263.4]
  wire [6:0] _T_88; // @[Counters.scala 47:33:freechips.rocketchip.system.DefaultRV32Config.fir@170263.4]
  reg [57:0] _T_89; // @[Counters.scala 51:27:freechips.rocketchip.system.DefaultRV32Config.fir@170265.4]
  reg [63:0] _RAND_84;
  wire  _T_90; // @[Counters.scala 52:20:freechips.rocketchip.system.DefaultRV32Config.fir@170266.4]
  wire [57:0] _T_92; // @[Counters.scala 52:43:freechips.rocketchip.system.DefaultRV32Config.fir@170269.6]
  wire [63:0] _T_93; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170272.4]
  wire  _T_94; // @[CSR.scala 403:103:freechips.rocketchip.system.DefaultRV32Config.fir@170273.4]
  reg [5:0] _T_95; // @[Counters.scala 46:37:freechips.rocketchip.system.DefaultRV32Config.fir@170274.4]
  reg [31:0] _RAND_85;
  wire [5:0] _GEN_441; // @[Counters.scala 47:33:freechips.rocketchip.system.DefaultRV32Config.fir@170275.4]
  wire [6:0] _T_96; // @[Counters.scala 47:33:freechips.rocketchip.system.DefaultRV32Config.fir@170275.4]
  reg [57:0] _T_97; // @[Counters.scala 51:27:freechips.rocketchip.system.DefaultRV32Config.fir@170277.4]
  reg [63:0] _RAND_86;
  wire  _T_98; // @[Counters.scala 52:20:freechips.rocketchip.system.DefaultRV32Config.fir@170278.4]
  wire [57:0] _T_100; // @[Counters.scala 52:43:freechips.rocketchip.system.DefaultRV32Config.fir@170281.6]
  wire [63:0] _T_101; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170284.4]
  wire [15:0] _T_116; // @[CSR.scala 416:22:freechips.rocketchip.system.DefaultRV32Config.fir@170306.4]
  wire [15:0] read_mip; // @[CSR.scala 416:29:freechips.rocketchip.system.DefaultRV32Config.fir@170307.4]
  wire [31:0] _GEN_442; // @[CSR.scala 419:56:freechips.rocketchip.system.DefaultRV32Config.fir@170308.4]
  wire [31:0] pending_interrupts; // @[CSR.scala 419:56:freechips.rocketchip.system.DefaultRV32Config.fir@170308.4]
  wire [14:0] d_interrupts; // @[CSR.scala 420:42:freechips.rocketchip.system.DefaultRV32Config.fir@170310.4]
  wire  _T_119; // @[CSR.scala 421:51:freechips.rocketchip.system.DefaultRV32Config.fir@170312.4]
  wire [31:0] _T_120; // @[CSR.scala 421:73:freechips.rocketchip.system.DefaultRV32Config.fir@170313.4]
  wire [31:0] _T_122; // @[CSR.scala 421:71:freechips.rocketchip.system.DefaultRV32Config.fir@170315.4]
  wire [31:0] m_interrupts; // @[CSR.scala 421:25:freechips.rocketchip.system.DefaultRV32Config.fir@170316.4]
  wire  _T_128; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170323.4]
  wire  _T_129; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170324.4]
  wire  _T_130; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170325.4]
  wire  _T_131; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170326.4]
  wire  _T_132; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170327.4]
  wire  _T_133; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170328.4]
  wire  _T_134; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170329.4]
  wire  _T_135; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170330.4]
  wire  _T_136; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170331.4]
  wire  _T_137; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170332.4]
  wire  _T_138; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170333.4]
  wire  _T_139; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170334.4]
  wire  _T_140; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170335.4]
  wire  _T_141; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170336.4]
  wire  _T_142; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170337.4]
  wire  _T_143; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170338.4]
  wire  _T_144; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170339.4]
  wire  _T_145; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170340.4]
  wire  _T_146; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170341.4]
  wire  _T_147; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170342.4]
  wire  _T_148; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170343.4]
  wire  _T_149; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170344.4]
  wire  _T_150; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170345.4]
  wire  _T_151; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170346.4]
  wire  _T_152; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170347.4]
  wire  _T_166; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170361.4]
  wire  _T_167; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170362.4]
  wire  _T_168; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170363.4]
  wire  _T_169; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170364.4]
  wire  _T_170; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170365.4]
  wire  _T_171; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170366.4]
  wire  _T_172; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170367.4]
  wire  _T_173; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170368.4]
  wire  _T_174; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170369.4]
  wire  _T_175; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170370.4]
  wire  _T_176; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170371.4]
  wire  _T_177; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170372.4]
  wire  _T_178; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170373.4]
  wire  _T_179; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170374.4]
  wire  _T_180; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170375.4]
  wire  _T_181; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170376.4]
  wire  _T_182; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170377.4]
  wire  _T_183; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170378.4]
  wire  _T_184; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170379.4]
  wire  _T_185; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170380.4]
  wire  _T_186; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170381.4]
  wire  _T_187; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170382.4]
  wire  _T_188; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170383.4]
  wire  anyInterrupt; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170384.4]
  wire [3:0] _T_253; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170449.4]
  wire [3:0] _T_254; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170450.4]
  wire [3:0] _T_255; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170451.4]
  wire [3:0] _T_256; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170452.4]
  wire [3:0] _T_257; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170453.4]
  wire [3:0] _T_258; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170454.4]
  wire [3:0] _T_259; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170455.4]
  wire [3:0] _T_260; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170456.4]
  wire [3:0] _T_261; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170457.4]
  wire [3:0] _T_262; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170458.4]
  wire [3:0] _T_263; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170459.4]
  wire [3:0] _T_264; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170460.4]
  wire [3:0] _T_265; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170461.4]
  wire [3:0] _T_266; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170462.4]
  wire [3:0] _T_267; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170463.4]
  wire [3:0] _T_268; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170464.4]
  wire [3:0] _T_269; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170465.4]
  wire [3:0] _T_270; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170466.4]
  wire [3:0] _T_271; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170467.4]
  wire [3:0] _T_272; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170468.4]
  wire [3:0] _T_273; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170469.4]
  wire [3:0] _T_274; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170470.4]
  wire [3:0] _T_275; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170471.4]
  wire [3:0] whichInterrupt; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170472.4]
  wire [31:0] _GEN_443; // @[CSR.scala 425:43:freechips.rocketchip.system.DefaultRV32Config.fir@170473.4]
  wire  _T_277; // @[CSR.scala 426:36:freechips.rocketchip.system.DefaultRV32Config.fir@170475.4]
  wire  _T_278; // @[CSR.scala 426:33:freechips.rocketchip.system.DefaultRV32Config.fir@170476.4]
  wire  _T_279; // @[CSR.scala 426:51:freechips.rocketchip.system.DefaultRV32Config.fir@170477.4]
  wire  _T_280; // @[CSR.scala 426:88:freechips.rocketchip.system.DefaultRV32Config.fir@170478.4]
  wire  _T_281; // @[CSR.scala 426:76:freechips.rocketchip.system.DefaultRV32Config.fir@170479.4]
  wire  _T_284; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170487.4]
  wire [30:0] _T_285; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170488.4]
  wire [30:0] _T_288; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170491.4]
  wire [30:0] _T_289; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170492.4]
  wire [30:0] _T_290; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170493.4]
  wire [32:0] _T_291; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170494.4]
  wire  _T_293; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170499.4]
  wire [30:0] _T_294; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170500.4]
  wire [30:0] _T_297; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170503.4]
  wire [30:0] _T_298; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170504.4]
  wire [30:0] _T_299; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170505.4]
  wire [32:0] _T_300; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170506.4]
  wire  _T_302; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170511.4]
  wire [30:0] _T_303; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170512.4]
  wire [30:0] _T_306; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170515.4]
  wire [30:0] _T_307; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170516.4]
  wire [30:0] _T_308; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170517.4]
  wire [32:0] _T_309; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170518.4]
  wire  _T_311; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170523.4]
  wire [30:0] _T_312; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170524.4]
  wire [30:0] _T_315; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170527.4]
  wire [30:0] _T_316; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170528.4]
  wire [30:0] _T_317; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170529.4]
  wire [32:0] _T_318; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170530.4]
  wire  _T_320; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170535.4]
  wire [30:0] _T_321; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170536.4]
  wire [30:0] _T_324; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170539.4]
  wire [30:0] _T_325; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170540.4]
  wire [30:0] _T_326; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170541.4]
  wire [32:0] _T_327; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170542.4]
  wire  _T_329; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170547.4]
  wire [30:0] _T_330; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170548.4]
  wire [30:0] _T_333; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170551.4]
  wire [30:0] _T_334; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170552.4]
  wire [30:0] _T_335; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170553.4]
  wire [32:0] _T_336; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170554.4]
  wire  _T_338; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170559.4]
  wire [30:0] _T_339; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170560.4]
  wire [30:0] _T_342; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170563.4]
  wire [30:0] _T_343; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170564.4]
  wire [30:0] _T_344; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170565.4]
  wire [32:0] _T_345; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170566.4]
  wire  _T_347; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170571.4]
  wire [30:0] _T_348; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170572.4]
  wire [30:0] _T_351; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170575.4]
  wire [30:0] _T_352; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170576.4]
  wire [30:0] _T_353; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170577.4]
  wire [32:0] _T_354; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170578.4]
  reg [31:0] reg_misa; // @[CSR.scala 444:21:freechips.rocketchip.system.DefaultRV32Config.fir@170588.4]
  reg [31:0] _RAND_87;
  wire [6:0] _T_360; // @[CSR.scala 445:38:freechips.rocketchip.system.DefaultRV32Config.fir@170594.4]
  wire [18:0] _T_368; // @[CSR.scala 445:38:freechips.rocketchip.system.DefaultRV32Config.fir@170602.4]
  wire [14:0] _T_375; // @[CSR.scala 445:38:freechips.rocketchip.system.DefaultRV32Config.fir@170609.4]
  wire [101:0] _T_384; // @[CSR.scala 445:38:freechips.rocketchip.system.DefaultRV32Config.fir@170618.4]
  wire [31:0] read_mstatus; // @[CSR.scala 445:40:freechips.rocketchip.system.DefaultRV32Config.fir@170619.4]
  wire  _T_385; // @[CSR.scala 1066:41:freechips.rocketchip.system.DefaultRV32Config.fir@170620.4]
  wire [6:0] _T_386; // @[CSR.scala 1066:39:freechips.rocketchip.system.DefaultRV32Config.fir@170621.4]
  wire [31:0] _T_388; // @[package.scala 131:41:freechips.rocketchip.system.DefaultRV32Config.fir@170623.4]
  wire [31:0] _T_389; // @[package.scala 131:37:freechips.rocketchip.system.DefaultRV32Config.fir@170624.4]
  wire [31:0] read_mtvec; // @[package.scala 131:35:freechips.rocketchip.system.DefaultRV32Config.fir@170625.4]
  wire [6:0] _T_400; // @[CSR.scala 451:48:freechips.rocketchip.system.DefaultRV32Config.fir@170637.4]
  wire [31:0] _T_408; // @[CSR.scala 451:48:freechips.rocketchip.system.DefaultRV32Config.fir@170645.4]
  wire [31:0] _T_409; // @[CSR.scala 1065:28:freechips.rocketchip.system.DefaultRV32Config.fir@170646.4]
  wire  _T_410; // @[CSR.scala 1065:45:freechips.rocketchip.system.DefaultRV32Config.fir@170647.4]
  wire [1:0] _T_411; // @[CSR.scala 1065:36:freechips.rocketchip.system.DefaultRV32Config.fir@170648.4]
  wire [31:0] _GEN_444; // @[CSR.scala 1065:31:freechips.rocketchip.system.DefaultRV32Config.fir@170649.4]
  wire [31:0] _T_412; // @[CSR.scala 1065:31:freechips.rocketchip.system.DefaultRV32Config.fir@170649.4]
  wire [31:0] _T_413; // @[CSR.scala 1065:26:freechips.rocketchip.system.DefaultRV32Config.fir@170650.4]
  wire [11:0] _T_419; // @[CSR.scala 465:27:freechips.rocketchip.system.DefaultRV32Config.fir@170656.4]
  wire [31:0] _T_426; // @[CSR.scala 465:27:freechips.rocketchip.system.DefaultRV32Config.fir@170663.4]
  wire [31:0] _T_427; // @[CSR.scala 1065:28:freechips.rocketchip.system.DefaultRV32Config.fir@170664.4]
  wire [31:0] _T_430; // @[CSR.scala 1065:31:freechips.rocketchip.system.DefaultRV32Config.fir@170667.4]
  wire [31:0] _T_431; // @[CSR.scala 1065:26:freechips.rocketchip.system.DefaultRV32Config.fir@170668.4]
  wire [7:0] _T_432; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170669.4]
  wire [8:0] _T_434; // @[CSR.scala 469:44:freechips.rocketchip.system.DefaultRV32Config.fir@170671.4]
  wire [9:0] read_fcsr; // @[CSR.scala 469:78:freechips.rocketchip.system.DefaultRV32Config.fir@170673.4]
  wire [31:0] _T_494; // @[CSR.scala 509:50:freechips.rocketchip.system.DefaultRV32Config.fir@170732.4]
  wire [31:0] _T_495; // @[CSR.scala 510:54:freechips.rocketchip.system.DefaultRV32Config.fir@170733.4]
  wire [7:0] _T_512; // @[package.scala 36:38:freechips.rocketchip.system.DefaultRV32Config.fir@170761.4]
  wire [7:0] _T_522; // @[package.scala 36:38:freechips.rocketchip.system.DefaultRV32Config.fir@170771.4]
  wire [15:0] _T_528; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170777.4]
  wire [31:0] _T_530; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170779.4]
  wire [7:0] _T_535; // @[package.scala 36:38:freechips.rocketchip.system.DefaultRV32Config.fir@170784.4]
  wire [7:0] _T_545; // @[package.scala 36:38:freechips.rocketchip.system.DefaultRV32Config.fir@170794.4]
  wire [15:0] _T_551; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170800.4]
  wire [31:0] _T_553; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170802.4]
  wire  _T_601; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170854.4]
  wire  _T_602; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170855.4]
  wire  _T_603; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170856.4]
  wire  _T_604; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170857.4]
  wire  _T_605; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170858.4]
  wire  _T_606; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170859.4]
  wire  _T_607; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170860.4]
  wire  _T_608; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170861.4]
  wire  _T_609; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170862.4]
  wire  _T_610; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170863.4]
  wire  _T_611; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170864.4]
  wire  _T_613; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170866.4]
  wire  _T_614; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170867.4]
  wire  _T_615; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170868.4]
  wire  _T_616; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170869.4]
  wire  _T_617; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170870.4]
  wire  _T_618; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170871.4]
  wire  _T_619; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170872.4]
  wire  _T_620; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170873.4]
  wire  _T_766; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171019.4]
  wire  _T_767; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171020.4]
  wire  _T_768; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171021.4]
  wire  _T_769; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171022.4]
  wire  _T_770; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171023.4]
  wire  _T_771; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171024.4]
  wire  _T_772; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171025.4]
  wire  _T_773; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171026.4]
  wire  _T_774; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171027.4]
  wire  _T_777; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171030.4]
  wire  _T_778; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171031.4]
  wire  _T_779; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171032.4]
  wire  _T_780; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171033.4]
  wire  _T_781; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171034.4]
  wire  _T_782; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171035.4]
  wire  _T_783; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171036.4]
  wire  _T_784; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171037.4]
  wire  _T_794; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171047.4]
  wire  _T_796; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171049.4]
  wire  _T_797; // @[CSR.scala 1043:13:freechips.rocketchip.system.DefaultRV32Config.fir@171050.4]
  wire [31:0] _T_798; // @[CSR.scala 1043:9:freechips.rocketchip.system.DefaultRV32Config.fir@171051.4]
  wire [31:0] _T_799; // @[CSR.scala 1043:34:freechips.rocketchip.system.DefaultRV32Config.fir@171052.4]
  wire [1:0] _T_800; // @[CSR.scala 1043:53:freechips.rocketchip.system.DefaultRV32Config.fir@171053.4]
  wire  _T_801; // @[CSR.scala 1043:59:freechips.rocketchip.system.DefaultRV32Config.fir@171054.4]
  wire [31:0] _T_802; // @[CSR.scala 1043:49:freechips.rocketchip.system.DefaultRV32Config.fir@171055.4]
  wire [31:0] _T_803; // @[CSR.scala 1043:45:freechips.rocketchip.system.DefaultRV32Config.fir@171056.4]
  wire [31:0] wdata; // @[CSR.scala 1043:43:freechips.rocketchip.system.DefaultRV32Config.fir@171057.4]
  wire [31:0] _T_814; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171069.4]
  wire  _T_815; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171070.4]
  wire [31:0] _T_817; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171072.4]
  wire  _T_818; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171073.4]
  wire  insn_cease; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171082.4]
  wire  insn_wfi; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171084.4]
  wire [31:0] _T_825; // @[CSR.scala 593:30:freechips.rocketchip.system.DefaultRV32Config.fir@171086.4]
  wire [31:0] _T_832; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171093.4]
  wire  _T_833; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171094.4]
  wire  _T_846; // @[CSR.scala 595:55:freechips.rocketchip.system.DefaultRV32Config.fir@171107.4]
  wire [4:0] _T_858; // @[CSR.scala 598:34:freechips.rocketchip.system.DefaultRV32Config.fir@171119.4]
  wire [31:0] _T_860; // @[CSR.scala 599:68:freechips.rocketchip.system.DefaultRV32Config.fir@171121.4]
  wire  _T_861; // @[CSR.scala 599:68:freechips.rocketchip.system.DefaultRV32Config.fir@171122.4]
  wire  _T_862; // @[CSR.scala 599:50:freechips.rocketchip.system.DefaultRV32Config.fir@171123.4]
  wire  _T_869; // @[CSR.scala 601:39:freechips.rocketchip.system.DefaultRV32Config.fir@171130.4]
  wire  _T_870; // @[CSR.scala 601:57:freechips.rocketchip.system.DefaultRV32Config.fir@171131.4]
  wire  _T_871; // @[CSR.scala 601:48:freechips.rocketchip.system.DefaultRV32Config.fir@171132.4]
  wire [11:0] _T_877; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171140.4]
  wire [1:0] _T_885; // @[CSR.scala 605:56:freechips.rocketchip.system.DefaultRV32Config.fir@171150.4]
  wire  _T_886; // @[CSR.scala 605:44:freechips.rocketchip.system.DefaultRV32Config.fir@171151.4]
  wire  _T_887; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171152.4]
  wire  _T_888; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171153.4]
  wire  _T_889; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171154.4]
  wire  _T_890; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171155.4]
  wire  _T_891; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171156.4]
  wire  _T_892; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171157.4]
  wire  _T_893; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171158.4]
  wire  _T_894; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171159.4]
  wire  _T_895; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171160.4]
  wire  _T_896; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171161.4]
  wire  _T_897; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171162.4]
  wire  _T_898; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171163.4]
  wire  _T_899; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171164.4]
  wire  _T_900; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171165.4]
  wire  _T_901; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171166.4]
  wire  _T_902; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171167.4]
  wire  _T_903; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171168.4]
  wire  _T_904; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171169.4]
  wire  _T_905; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171170.4]
  wire  _T_906; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171171.4]
  wire  _T_907; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171172.4]
  wire  _T_908; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171173.4]
  wire  _T_909; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171174.4]
  wire  _T_910; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171175.4]
  wire  _T_911; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171176.4]
  wire  _T_912; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171177.4]
  wire  _T_913; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171178.4]
  wire  _T_914; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171179.4]
  wire  _T_915; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171180.4]
  wire  _T_916; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171181.4]
  wire  _T_917; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171182.4]
  wire  _T_918; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171183.4]
  wire  _T_919; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171184.4]
  wire  _T_920; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171185.4]
  wire  _T_921; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171186.4]
  wire  _T_922; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171187.4]
  wire  _T_923; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171188.4]
  wire  _T_924; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171189.4]
  wire  _T_925; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171190.4]
  wire  _T_926; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171191.4]
  wire  _T_927; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171192.4]
  wire  _T_928; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171193.4]
  wire  _T_929; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171194.4]
  wire  _T_930; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171195.4]
  wire  _T_931; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171196.4]
  wire  _T_932; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171197.4]
  wire  _T_933; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171198.4]
  wire  _T_934; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171199.4]
  wire  _T_935; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171200.4]
  wire  _T_936; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171201.4]
  wire  _T_937; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171202.4]
  wire  _T_938; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171203.4]
  wire  _T_939; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171204.4]
  wire  _T_940; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171205.4]
  wire  _T_941; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171206.4]
  wire  _T_942; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171207.4]
  wire  _T_943; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171208.4]
  wire  _T_944; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171209.4]
  wire  _T_945; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171210.4]
  wire  _T_946; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171211.4]
  wire  _T_947; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171212.4]
  wire  _T_948; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171213.4]
  wire  _T_949; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171214.4]
  wire  _T_950; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171215.4]
  wire  _T_951; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171216.4]
  wire  _T_952; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171217.4]
  wire  _T_953; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171218.4]
  wire  _T_954; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171219.4]
  wire  _T_955; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171220.4]
  wire  _T_956; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171221.4]
  wire  _T_957; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171222.4]
  wire  _T_958; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171223.4]
  wire  _T_959; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171224.4]
  wire  _T_960; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171225.4]
  wire  _T_961; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171226.4]
  wire  _T_962; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171227.4]
  wire  _T_963; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171228.4]
  wire  _T_964; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171229.4]
  wire  _T_965; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171230.4]
  wire  _T_966; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171231.4]
  wire  _T_967; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171232.4]
  wire  _T_968; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171233.4]
  wire  _T_969; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171234.4]
  wire  _T_970; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171235.4]
  wire  _T_971; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171236.4]
  wire  _T_972; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171237.4]
  wire  _T_973; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171238.4]
  wire  _T_974; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171239.4]
  wire  _T_975; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171240.4]
  wire  _T_976; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171241.4]
  wire  _T_977; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171242.4]
  wire  _T_978; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171243.4]
  wire  _T_979; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171244.4]
  wire  _T_980; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171245.4]
  wire  _T_981; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171246.4]
  wire  _T_982; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171247.4]
  wire  _T_983; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171248.4]
  wire  _T_984; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171249.4]
  wire  _T_985; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171250.4]
  wire  _T_986; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171251.4]
  wire  _T_987; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171252.4]
  wire  _T_988; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171253.4]
  wire  _T_989; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171254.4]
  wire  _T_990; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171255.4]
  wire  _T_991; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171256.4]
  wire  _T_992; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171257.4]
  wire  _T_993; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171258.4]
  wire  _T_994; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171259.4]
  wire  _T_995; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171260.4]
  wire  _T_996; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171261.4]
  wire  _T_997; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171262.4]
  wire  _T_998; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171263.4]
  wire  _T_999; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171264.4]
  wire  _T_1000; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171265.4]
  wire  _T_1001; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171266.4]
  wire  _T_1002; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171267.4]
  wire  _T_1003; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171268.4]
  wire  _T_1004; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171269.4]
  wire  _T_1005; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171270.4]
  wire  _T_1006; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171271.4]
  wire  _T_1007; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171272.4]
  wire  _T_1008; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171273.4]
  wire  _T_1009; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171274.4]
  wire  _T_1010; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171275.4]
  wire  _T_1011; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171276.4]
  wire  _T_1012; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171277.4]
  wire  _T_1013; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171278.4]
  wire  _T_1014; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171279.4]
  wire  _T_1015; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171280.4]
  wire  _T_1016; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171281.4]
  wire  _T_1017; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171282.4]
  wire  _T_1018; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171283.4]
  wire  _T_1019; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171284.4]
  wire  _T_1020; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171285.4]
  wire  _T_1021; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171286.4]
  wire  _T_1022; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171287.4]
  wire  _T_1023; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171288.4]
  wire  _T_1024; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171289.4]
  wire  _T_1025; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171290.4]
  wire  _T_1026; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171291.4]
  wire  _T_1027; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171292.4]
  wire  _T_1028; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171293.4]
  wire  _T_1029; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171294.4]
  wire  _T_1030; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171295.4]
  wire  _T_1031; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171296.4]
  wire  _T_1032; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171297.4]
  wire  _T_1033; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171298.4]
  wire  _T_1034; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171299.4]
  wire  _T_1035; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171300.4]
  wire  _T_1036; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171301.4]
  wire  _T_1037; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171302.4]
  wire  _T_1038; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171303.4]
  wire  _T_1039; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171304.4]
  wire  _T_1040; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171305.4]
  wire  _T_1041; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171306.4]
  wire  _T_1042; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171307.4]
  wire  _T_1043; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171308.4]
  wire  _T_1044; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171309.4]
  wire  _T_1045; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171310.4]
  wire  _T_1046; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171311.4]
  wire  _T_1047; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171312.4]
  wire  _T_1048; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171313.4]
  wire  _T_1049; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171314.4]
  wire  _T_1050; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171315.4]
  wire  _T_1051; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171316.4]
  wire  _T_1052; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171317.4]
  wire  _T_1053; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171318.4]
  wire  _T_1054; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171319.4]
  wire  _T_1055; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171320.4]
  wire  _T_1056; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171321.4]
  wire  _T_1057; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171322.4]
  wire  _T_1058; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171323.4]
  wire  _T_1059; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171324.4]
  wire  _T_1060; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171325.4]
  wire  _T_1061; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171326.4]
  wire  _T_1062; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171327.4]
  wire  _T_1063; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171328.4]
  wire  _T_1064; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171329.4]
  wire  _T_1065; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171330.4]
  wire  _T_1066; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171331.4]
  wire  _T_1067; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171332.4]
  wire  _T_1068; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171333.4]
  wire  _T_1069; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171334.4]
  wire  _T_1070; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171335.4]
  wire  _T_1071; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171336.4]
  wire  _T_1072; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171337.4]
  wire  _T_1073; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171338.4]
  wire  _T_1074; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171339.4]
  wire  _T_1075; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171340.4]
  wire  _T_1076; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171341.4]
  wire  _T_1077; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171342.4]
  wire  _T_1078; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171343.4]
  wire  _T_1079; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171344.4]
  wire  _T_1080; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171345.4]
  wire  _T_1081; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171346.4]
  wire  _T_1082; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171347.4]
  wire  _T_1083; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171348.4]
  wire  _T_1084; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171349.4]
  wire  _T_1085; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171350.4]
  wire  _T_1086; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171351.4]
  wire  _T_1087; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171352.4]
  wire  _T_1088; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171353.4]
  wire  _T_1089; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171354.4]
  wire  _T_1090; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171355.4]
  wire  _T_1091; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171356.4]
  wire  _T_1092; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171357.4]
  wire  _T_1093; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171358.4]
  wire  _T_1094; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171359.4]
  wire  _T_1095; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171360.4]
  wire  _T_1096; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171361.4]
  wire  _T_1097; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171362.4]
  wire  _T_1098; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171363.4]
  wire  _T_1099; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171364.4]
  wire  _T_1100; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171365.4]
  wire  _T_1101; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171366.4]
  wire  _T_1102; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171367.4]
  wire  _T_1103; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171368.4]
  wire  _T_1104; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171369.4]
  wire  _T_1105; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171370.4]
  wire  _T_1106; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171371.4]
  wire  _T_1107; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171372.4]
  wire  _T_1108; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171373.4]
  wire  _T_1109; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171374.4]
  wire  _T_1110; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171375.4]
  wire  _T_1111; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171376.4]
  wire  _T_1112; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171377.4]
  wire  _T_1113; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171378.4]
  wire  _T_1114; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171379.4]
  wire  _T_1115; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171380.4]
  wire  _T_1116; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171381.4]
  wire  _T_1117; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171382.4]
  wire  _T_1118; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171383.4]
  wire  _T_1119; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171384.4]
  wire  _T_1120; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171385.4]
  wire  _T_1121; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171386.4]
  wire  _T_1122; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171387.4]
  wire  _T_1123; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171388.4]
  wire  _T_1124; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171389.4]
  wire  _T_1125; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171390.4]
  wire  _T_1126; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171391.4]
  wire  _T_1127; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171392.4]
  wire  _T_1128; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171393.4]
  wire  _T_1129; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171394.4]
  wire  _T_1130; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171395.4]
  wire  _T_1131; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171396.4]
  wire  _T_1132; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171397.4]
  wire  _T_1133; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171398.4]
  wire  _T_1134; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171399.4]
  wire  _T_1135; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171400.4]
  wire  _T_1136; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171401.4]
  wire  _T_1137; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171402.4]
  wire  _T_1138; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171403.4]
  wire  _T_1139; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171404.4]
  wire  _T_1140; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171405.4]
  wire  _T_1141; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171406.4]
  wire  _T_1142; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171407.4]
  wire  _T_1143; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171408.4]
  wire  _T_1144; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171409.4]
  wire  _T_1145; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171410.4]
  wire  _T_1146; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171411.4]
  wire  _T_1147; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171412.4]
  wire  _T_1148; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171413.4]
  wire  _T_1149; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171414.4]
  wire  _T_1150; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171415.4]
  wire  _T_1151; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171416.4]
  wire  _T_1152; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171417.4]
  wire  _T_1153; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171418.4]
  wire  _T_1154; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171419.4]
  wire  _T_1155; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171420.4]
  wire  _T_1156; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171421.4]
  wire  _T_1157; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171422.4]
  wire  _T_1158; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171423.4]
  wire  _T_1159; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171424.4]
  wire  _T_1160; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171425.4]
  wire  _T_1161; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171426.4]
  wire  _T_1162; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171427.4]
  wire  _T_1163; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171428.4]
  wire  _T_1164; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171429.4]
  wire  _T_1165; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171430.4]
  wire  _T_1166; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171431.4]
  wire  _T_1167; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171432.4]
  wire  _T_1168; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171433.4]
  wire  _T_1169; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171434.4]
  wire  _T_1170; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171435.4]
  wire  _T_1171; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171436.4]
  wire  _T_1172; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171437.4]
  wire  _T_1173; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171438.4]
  wire  _T_1174; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171439.4]
  wire  _T_1175; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171440.4]
  wire  _T_1176; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171441.4]
  wire  _T_1177; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171442.4]
  wire  _T_1178; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171443.4]
  wire  _T_1179; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171444.4]
  wire  _T_1180; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171445.4]
  wire  _T_1181; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171446.4]
  wire  _T_1182; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171447.4]
  wire  _T_1183; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171448.4]
  wire  _T_1184; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171449.4]
  wire  _T_1185; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171450.4]
  wire  _T_1186; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171451.4]
  wire  _T_1187; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171452.4]
  wire  _T_1188; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171453.4]
  wire  _T_1189; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171454.4]
  wire  _T_1190; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171455.4]
  wire  _T_1191; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171456.4]
  wire  _T_1192; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171457.4]
  wire  _T_1193; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171458.4]
  wire  _T_1194; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171459.4]
  wire  _T_1195; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171460.4]
  wire  _T_1196; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171461.4]
  wire  _T_1197; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171462.4]
  wire  _T_1198; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171463.4]
  wire  _T_1199; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171464.4]
  wire  _T_1200; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171465.4]
  wire  _T_1201; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171466.4]
  wire  _T_1202; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171467.4]
  wire  _T_1203; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171468.4]
  wire  _T_1204; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171469.4]
  wire  _T_1205; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171470.4]
  wire  _T_1206; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171471.4]
  wire  _T_1207; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171472.4]
  wire  _T_1208; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171473.4]
  wire  _T_1209; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171474.4]
  wire  _T_1210; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171475.4]
  wire  _T_1211; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171476.4]
  wire  _T_1212; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171477.4]
  wire  _T_1213; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171478.4]
  wire  _T_1214; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171479.4]
  wire  _T_1215; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171480.4]
  wire  _T_1216; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171481.4]
  wire  _T_1217; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171482.4]
  wire  _T_1218; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171483.4]
  wire  _T_1219; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171484.4]
  wire  _T_1220; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171485.4]
  wire  _T_1221; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171486.4]
  wire  _T_1222; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171487.4]
  wire  _T_1223; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171488.4]
  wire  _T_1224; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171489.4]
  wire  _T_1225; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171490.4]
  wire  _T_1226; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171491.4]
  wire  _T_1227; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171492.4]
  wire  _T_1228; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171493.4]
  wire  _T_1229; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171494.4]
  wire  _T_1230; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171495.4]
  wire  _T_1231; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171496.4]
  wire  _T_1232; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171497.4]
  wire  _T_1233; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171498.4]
  wire  _T_1234; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171499.4]
  wire  _T_1235; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171500.4]
  wire  _T_1236; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171501.4]
  wire  _T_1237; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171502.4]
  wire  _T_1238; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171503.4]
  wire  _T_1239; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171504.4]
  wire  _T_1240; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171505.4]
  wire  _T_1241; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171506.4]
  wire  _T_1242; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171507.4]
  wire  _T_1243; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171508.4]
  wire  _T_1244; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171509.4]
  wire  _T_1245; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171510.4]
  wire  _T_1246; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171511.4]
  wire  _T_1247; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171512.4]
  wire  _T_1248; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171513.4]
  wire  _T_1249; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171514.4]
  wire  _T_1250; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171515.4]
  wire  _T_1251; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171516.4]
  wire  _T_1252; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171517.4]
  wire  _T_1253; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171518.4]
  wire  _T_1254; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171519.4]
  wire  _T_1255; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171520.4]
  wire  _T_1256; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171521.4]
  wire  _T_1257; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171522.4]
  wire  _T_1258; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171523.4]
  wire  _T_1259; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171524.4]
  wire  _T_1260; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171525.4]
  wire  _T_1261; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171526.4]
  wire  _T_1262; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171527.4]
  wire  _T_1263; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171528.4]
  wire  _T_1264; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171529.4]
  wire  _T_1265; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171530.4]
  wire  _T_1266; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171531.4]
  wire  _T_1267; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171532.4]
  wire  _T_1268; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171533.4]
  wire  _T_1269; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171534.4]
  wire  _T_1270; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171535.4]
  wire  _T_1271; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171536.4]
  wire  _T_1272; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171537.4]
  wire  _T_1273; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171538.4]
  wire  _T_1274; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171539.4]
  wire  _T_1275; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171540.4]
  wire  _T_1276; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171541.4]
  wire  _T_1277; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171542.4]
  wire  _T_1278; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171543.4]
  wire  _T_1279; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171544.4]
  wire  _T_1280; // @[CSR.scala 606:7:freechips.rocketchip.system.DefaultRV32Config.fir@171545.4]
  wire  _T_1281; // @[CSR.scala 605:62:freechips.rocketchip.system.DefaultRV32Config.fir@171546.4]
  wire  _T_1286; // @[package.scala 162:47:freechips.rocketchip.system.DefaultRV32Config.fir@171551.4]
  wire  _T_1287; // @[package.scala 162:60:freechips.rocketchip.system.DefaultRV32Config.fir@171552.4]
  wire  _T_1288; // @[package.scala 162:55:freechips.rocketchip.system.DefaultRV32Config.fir@171553.4]
  wire  _T_1289; // @[package.scala 162:47:freechips.rocketchip.system.DefaultRV32Config.fir@171554.4]
  wire  _T_1290; // @[package.scala 162:60:freechips.rocketchip.system.DefaultRV32Config.fir@171555.4]
  wire  _T_1291; // @[package.scala 162:55:freechips.rocketchip.system.DefaultRV32Config.fir@171556.4]
  wire  _T_1292; // @[CSR.scala 608:66:freechips.rocketchip.system.DefaultRV32Config.fir@171557.4]
  wire  _T_1293; // @[CSR.scala 608:133:freechips.rocketchip.system.DefaultRV32Config.fir@171558.4]
  wire  _T_1294; // @[CSR.scala 608:130:freechips.rocketchip.system.DefaultRV32Config.fir@171559.4]
  wire  _T_1295; // @[CSR.scala 607:53:freechips.rocketchip.system.DefaultRV32Config.fir@171560.4]
  wire [11:0] _T_1296; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171561.4]
  wire  _T_1297; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171562.4]
  wire  _T_1301; // @[CSR.scala 609:42:freechips.rocketchip.system.DefaultRV32Config.fir@171566.4]
  wire  _T_1302; // @[CSR.scala 608:148:freechips.rocketchip.system.DefaultRV32Config.fir@171567.4]
  wire  _T_1305; // @[CSR.scala 611:21:freechips.rocketchip.system.DefaultRV32Config.fir@171570.4]
  wire [1:0] _T_1307; // @[CSR.scala 612:39:freechips.rocketchip.system.DefaultRV32Config.fir@171573.4]
  wire  _T_1309; // @[CSR.scala 613:40:freechips.rocketchip.system.DefaultRV32Config.fir@171576.4]
  wire  _T_1310; // @[CSR.scala 613:71:freechips.rocketchip.system.DefaultRV32Config.fir@171577.4]
  wire  _T_1311; // @[CSR.scala 613:57:freechips.rocketchip.system.DefaultRV32Config.fir@171578.4]
  wire  _T_1312; // @[CSR.scala 613:99:freechips.rocketchip.system.DefaultRV32Config.fir@171579.4]
  wire  _T_1313; // @[CSR.scala 613:130:freechips.rocketchip.system.DefaultRV32Config.fir@171580.4]
  wire  _T_1314; // @[CSR.scala 613:116:freechips.rocketchip.system.DefaultRV32Config.fir@171581.4]
  wire  _T_1315; // @[CSR.scala 613:85:freechips.rocketchip.system.DefaultRV32Config.fir@171582.4]
  wire  _T_1325; // @[CSR.scala 617:27:freechips.rocketchip.system.DefaultRV32Config.fir@171593.4]
  wire  _T_1326; // @[CSR.scala 617:14:freechips.rocketchip.system.DefaultRV32Config.fir@171594.4]
  wire  _T_1328; // @[CSR.scala 617:32:freechips.rocketchip.system.DefaultRV32Config.fir@171596.4]
  wire [11:0] _T_1353; // @[CSR.scala 629:37:freechips.rocketchip.system.DefaultRV32Config.fir@171628.4]
  wire [11:0] debugTVec; // @[CSR.scala 629:22:freechips.rocketchip.system.DefaultRV32Config.fir@171629.4]
  wire [4:0] _T_1363; // @[CSR.scala 638:32:freechips.rocketchip.system.DefaultRV32Config.fir@171640.4]
  wire [6:0] _T_1364; // @[CSR.scala 638:59:freechips.rocketchip.system.DefaultRV32Config.fir@171641.4]
  wire [24:0] _T_1365; // @[CSR.scala 639:33:freechips.rocketchip.system.DefaultRV32Config.fir@171642.4]
  wire [31:0] _T_1366; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@171643.4]
  wire  _T_1367; // @[CSR.scala 640:24:freechips.rocketchip.system.DefaultRV32Config.fir@171644.4]
  wire  _T_1369; // @[CSR.scala 640:28:freechips.rocketchip.system.DefaultRV32Config.fir@171646.4]
  wire [2:0] _T_1370; // @[CSR.scala 640:70:freechips.rocketchip.system.DefaultRV32Config.fir@171647.4]
  wire  _T_1371; // @[CSR.scala 640:94:freechips.rocketchip.system.DefaultRV32Config.fir@171648.4]
  wire  _T_1372; // @[CSR.scala 640:55:freechips.rocketchip.system.DefaultRV32Config.fir@171649.4]
  wire [29:0] _T_1373; // @[CSR.scala 641:38:freechips.rocketchip.system.DefaultRV32Config.fir@171650.4]
  wire [31:0] _T_1374; // @[CSR.scala 641:56:freechips.rocketchip.system.DefaultRV32Config.fir@171651.4]
  wire [31:0] notDebugTVec; // @[CSR.scala 641:8:freechips.rocketchip.system.DefaultRV32Config.fir@171652.4]
  wire [31:0] tvec; // @[CSR.scala 643:17:freechips.rocketchip.system.DefaultRV32Config.fir@171653.4]
  wire  _T_1379; // @[CSR.scala 649:32:freechips.rocketchip.system.DefaultRV32Config.fir@171663.4]
  wire  _T_1380; // @[CSR.scala 649:53:freechips.rocketchip.system.DefaultRV32Config.fir@171664.4]
  wire  _T_1381; // @[CSR.scala 649:37:freechips.rocketchip.system.DefaultRV32Config.fir@171665.4]
  wire  _T_1382; // @[CSR.scala 649:74:freechips.rocketchip.system.DefaultRV32Config.fir@171666.4]
  wire  _T_1385; // @[CSR.scala 654:53:freechips.rocketchip.system.DefaultRV32Config.fir@171674.4]
  reg [1:0] _T_1387; // @[CSR.scala 654:24:freechips.rocketchip.system.DefaultRV32Config.fir@171676.4]
  reg [31:0] _RAND_88;
  wire [1:0] _T_1389; // @[Bitwise.scala 47:55:freechips.rocketchip.system.DefaultRV32Config.fir@171682.4]
  wire [1:0] _T_1391; // @[Bitwise.scala 47:55:freechips.rocketchip.system.DefaultRV32Config.fir@171684.4]
  wire [2:0] _T_1393; // @[Bitwise.scala 47:55:freechips.rocketchip.system.DefaultRV32Config.fir@171686.4]
  wire  _T_1395; // @[CSR.scala 659:79:freechips.rocketchip.system.DefaultRV32Config.fir@171688.4]
  wire  _T_1397; // @[CSR.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@171690.4]
  wire  _T_1398; // @[CSR.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@171691.4]
  wire  _T_1400; // @[CSR.scala 661:18:freechips.rocketchip.system.DefaultRV32Config.fir@171697.4]
  wire  _T_1402; // @[CSR.scala 661:36:freechips.rocketchip.system.DefaultRV32Config.fir@171699.4]
  wire  _GEN_34; // @[CSR.scala 661:51:freechips.rocketchip.system.DefaultRV32Config.fir@171700.4]
  wire  _T_1403; // @[CSR.scala 662:28:freechips.rocketchip.system.DefaultRV32Config.fir@171703.4]
  wire  _T_1404; // @[CSR.scala 662:32:freechips.rocketchip.system.DefaultRV32Config.fir@171704.4]
  wire  _T_1405; // @[CSR.scala 662:55:freechips.rocketchip.system.DefaultRV32Config.fir@171705.4]
  wire  _T_1407; // @[CSR.scala 664:22:freechips.rocketchip.system.DefaultRV32Config.fir@171710.4]
  wire  _GEN_36; // @[CSR.scala 664:36:freechips.rocketchip.system.DefaultRV32Config.fir@171711.4]
  wire  _T_1415; // @[CSR.scala 667:10:freechips.rocketchip.system.DefaultRV32Config.fir@171728.4]
  wire  _T_1416; // @[CSR.scala 667:42:freechips.rocketchip.system.DefaultRV32Config.fir@171729.4]
  wire  _T_1417; // @[CSR.scala 667:29:freechips.rocketchip.system.DefaultRV32Config.fir@171730.4]
  wire  _T_1419; // @[CSR.scala 667:9:freechips.rocketchip.system.DefaultRV32Config.fir@171732.4]
  wire  _T_1420; // @[CSR.scala 667:9:freechips.rocketchip.system.DefaultRV32Config.fir@171733.4]
  wire [31:0] _T_1421; // @[CSR.scala 1064:28:freechips.rocketchip.system.DefaultRV32Config.fir@171738.4]
  wire [31:0] _T_1422; // @[CSR.scala 1064:31:freechips.rocketchip.system.DefaultRV32Config.fir@171739.4]
  wire [31:0] epc; // @[CSR.scala 1064:26:freechips.rocketchip.system.DefaultRV32Config.fir@171740.4]
  wire [1:0] _T_1424; // @[CSR.scala 678:86:freechips.rocketchip.system.DefaultRV32Config.fir@171750.10]
  wire [1:0] _T_1425; // @[CSR.scala 678:56:freechips.rocketchip.system.DefaultRV32Config.fir@171751.10]
  wire  _T_1427; // @[CSR.scala 1048:37:freechips.rocketchip.system.DefaultRV32Config.fir@171754.10]
  wire [1:0] _T_1429; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@171756.10]
  wire  _GEN_38; // @[CSR.scala 675:25:freechips.rocketchip.system.DefaultRV32Config.fir@171747.8]
  wire [1:0] _GEN_48; // @[CSR.scala 682:27:freechips.rocketchip.system.DefaultRV32Config.fir@171762.8]
  wire [1:0] _GEN_67; // @[CSR.scala 674:24:freechips.rocketchip.system.DefaultRV32Config.fir@171745.6]
  wire  _GEN_74; // @[CSR.scala 674:24:freechips.rocketchip.system.DefaultRV32Config.fir@171745.6]
  wire [1:0] _GEN_85; // @[CSR.scala 673:20:freechips.rocketchip.system.DefaultRV32Config.fir@171744.4]
  wire [31:0] _GEN_95; // @[CSR.scala 729:53:freechips.rocketchip.system.DefaultRV32Config.fir@172093.8]
  reg  _T_1743; // @[Reg.scala 27:20:freechips.rocketchip.system.DefaultRV32Config.fir@172120.4]
  reg [31:0] _RAND_89;
  wire  _GEN_117; // @[Reg.scala 28:19:freechips.rocketchip.system.DefaultRV32Config.fir@172121.4]
  wire [31:0] _T_1745; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172138.4]
  wire [31:0] _T_1746; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172139.4]
  wire [31:0] _T_1747; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172140.4]
  wire [31:0] _T_1748; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172141.4]
  wire [31:0] _T_1749; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172142.4]
  wire [15:0] _T_1750; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172143.4]
  wire [31:0] _T_1751; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172144.4]
  wire [31:0] _T_1752; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172145.4]
  wire [31:0] _T_1753; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172146.4]
  wire [31:0] _T_1754; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172147.4]
  wire [31:0] _T_1755; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172148.4]
  wire [31:0] _T_1757; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172150.4]
  wire [31:0] _T_1758; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172151.4]
  wire [31:0] _T_1759; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172152.4]
  wire [4:0] _T_1760; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172153.4]
  wire [2:0] _T_1761; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172154.4]
  wire [9:0] _T_1762; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172155.4]
  wire [63:0] _T_1763; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172156.4]
  wire [63:0] _T_1764; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172157.4]
  wire [31:0] _T_1910; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172303.4]
  wire [63:0] _T_1911; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172304.4]
  wire [63:0] _T_1912; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172305.4]
  wire [31:0] _T_1913; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172306.4]
  wire [31:0] _T_1914; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172307.4]
  wire [31:0] _T_1915; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172308.4]
  wire [31:0] _T_1916; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172309.4]
  wire [31:0] _T_1917; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172310.4]
  wire [31:0] _T_1918; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172311.4]
  wire [29:0] _T_1921; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172314.4]
  wire [29:0] _T_1922; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172315.4]
  wire [29:0] _T_1923; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172316.4]
  wire [29:0] _T_1924; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172317.4]
  wire [29:0] _T_1925; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172318.4]
  wire [29:0] _T_1926; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172319.4]
  wire [29:0] _T_1927; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172320.4]
  wire [29:0] _T_1928; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172321.4]
  wire [31:0] _T_1938; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172331.4]
  wire [31:0] _T_1940; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172333.4]
  wire [31:0] _T_1942; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172335.4]
  wire [31:0] _T_1943; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172336.4]
  wire [31:0] _T_1944; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172337.4]
  wire [31:0] _T_1945; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172338.4]
  wire [31:0] _GEN_448; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172339.4]
  wire [31:0] _T_1946; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172339.4]
  wire [31:0] _T_1947; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172340.4]
  wire [31:0] _T_1948; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172341.4]
  wire [31:0] _T_1949; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172342.4]
  wire [31:0] _T_1950; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172343.4]
  wire [31:0] _T_1951; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172344.4]
  wire [31:0] _T_1953; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172346.4]
  wire [31:0] _T_1954; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172347.4]
  wire [31:0] _T_1955; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172348.4]
  wire [31:0] _GEN_449; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172349.4]
  wire [31:0] _T_1956; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172349.4]
  wire [31:0] _GEN_450; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172350.4]
  wire [31:0] _T_1957; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172350.4]
  wire [31:0] _GEN_451; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172351.4]
  wire [31:0] _T_1958; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172351.4]
  wire [63:0] _GEN_452; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172352.4]
  wire [63:0] _T_1959; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172352.4]
  wire [63:0] _T_1960; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172353.4]
  wire [63:0] _GEN_453; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172499.4]
  wire [63:0] _T_2106; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172499.4]
  wire [63:0] _T_2107; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172500.4]
  wire [63:0] _T_2108; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172501.4]
  wire [63:0] _GEN_454; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172502.4]
  wire [63:0] _T_2109; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172502.4]
  wire [63:0] _GEN_455; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172503.4]
  wire [63:0] _T_2110; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172503.4]
  wire [63:0] _GEN_456; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172504.4]
  wire [63:0] _T_2111; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172504.4]
  wire [63:0] _GEN_457; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172505.4]
  wire [63:0] _T_2112; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172505.4]
  wire [63:0] _GEN_458; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172506.4]
  wire [63:0] _T_2113; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172506.4]
  wire [63:0] _GEN_459; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172507.4]
  wire [63:0] _T_2114; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172507.4]
  wire [63:0] _GEN_460; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172510.4]
  wire [63:0] _T_2117; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172510.4]
  wire [63:0] _GEN_461; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172511.4]
  wire [63:0] _T_2118; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172511.4]
  wire [63:0] _GEN_462; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172512.4]
  wire [63:0] _T_2119; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172512.4]
  wire [63:0] _GEN_463; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172513.4]
  wire [63:0] _T_2120; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172513.4]
  wire [63:0] _GEN_464; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172514.4]
  wire [63:0] _T_2121; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172514.4]
  wire [63:0] _GEN_465; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172515.4]
  wire [63:0] _T_2122; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172515.4]
  wire [63:0] _GEN_466; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172516.4]
  wire [63:0] _T_2123; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172516.4]
  wire [63:0] _GEN_467; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172517.4]
  wire [63:0] _T_2124; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172517.4]
  wire [63:0] _GEN_468; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172527.4]
  wire [63:0] _T_2134; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172527.4]
  wire [63:0] _GEN_469; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172529.4]
  wire [63:0] _T_2136; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172529.4]
  wire  _T_2140; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@172536.6]
  wire  _T_2141; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@172537.6]
  wire  _T_2142; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@172538.6]
  wire [4:0] _T_4502; // @[CSR.scala 781:30:freechips.rocketchip.system.DefaultRV32Config.fir@175693.6]
  wire [4:0] _GEN_118; // @[CSR.scala 780:30:freechips.rocketchip.system.DefaultRV32Config.fir@175692.4]
  wire  _T_4506; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@175700.4]
  wire  csr_wen; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@175701.4]
  wire [101:0] _T_4520; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175719.8 :freechips.rocketchip.system.DefaultRV32Config.fir@175721.8]
  wire  _T_4524; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175728.8]
  wire  _T_4528; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175736.8]
  wire [1:0] _T_4531; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175742.8]
  wire [1:0] _T_4532; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175744.8]
  wire  _T_4534; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175748.8]
  wire  _T_4552; // @[CSR.scala 1048:37:freechips.rocketchip.system.DefaultRV32Config.fir@175787.8]
  wire  _T_4555; // @[CSR.scala 1068:73:freechips.rocketchip.system.DefaultRV32Config.fir@175791.8]
  wire  _T_4558; // @[CSR.scala 821:20:freechips.rocketchip.system.DefaultRV32Config.fir@175798.8]
  wire  _T_4559; // @[CSR.scala 823:39:freechips.rocketchip.system.DefaultRV32Config.fir@175799.8]
  wire  _T_4560; // @[CSR.scala 823:33:freechips.rocketchip.system.DefaultRV32Config.fir@175800.8]
  wire  _T_4562; // @[CSR.scala 823:51:freechips.rocketchip.system.DefaultRV32Config.fir@175802.8]
  wire  _T_4563; // @[CSR.scala 823:43:freechips.rocketchip.system.DefaultRV32Config.fir@175803.8]
  wire [31:0] _T_4564; // @[CSR.scala 825:25:freechips.rocketchip.system.DefaultRV32Config.fir@175805.10]
  wire  _T_4565; // @[CSR.scala 825:35:freechips.rocketchip.system.DefaultRV32Config.fir@175806.10]
  wire [3:0] _T_4566; // @[CSR.scala 825:38:freechips.rocketchip.system.DefaultRV32Config.fir@175807.10]
  wire [31:0] _GEN_470; // @[CSR.scala 825:32:freechips.rocketchip.system.DefaultRV32Config.fir@175808.10]
  wire [31:0] _T_4567; // @[CSR.scala 825:32:freechips.rocketchip.system.DefaultRV32Config.fir@175808.10]
  wire [31:0] _T_4568; // @[CSR.scala 825:23:freechips.rocketchip.system.DefaultRV32Config.fir@175809.10]
  wire [31:0] _T_4569; // @[CSR.scala 825:55:freechips.rocketchip.system.DefaultRV32Config.fir@175810.10]
  wire [31:0] _T_4571; // @[CSR.scala 825:73:freechips.rocketchip.system.DefaultRV32Config.fir@175812.10]
  wire [31:0] _T_4572; // @[CSR.scala 825:62:freechips.rocketchip.system.DefaultRV32Config.fir@175813.10]
  wire [31:0] _T_4614; // @[CSR.scala 840:59:freechips.rocketchip.system.DefaultRV32Config.fir@175880.8]
  wire [31:0] _T_4616; // @[CSR.scala 1064:31:freechips.rocketchip.system.DefaultRV32Config.fir@175885.8]
  wire [31:0] _T_4617; // @[CSR.scala 1064:26:freechips.rocketchip.system.DefaultRV32Config.fir@175886.8]
  wire [31:0] _T_4618; // @[CSR.scala 845:62:freechips.rocketchip.system.DefaultRV32Config.fir@175896.8]
  wire [31:0] _T_4620; // @[CSR.scala 1058:47:freechips.rocketchip.system.DefaultRV32Config.fir@175904.8]
  wire [63:0] _T_4621; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@175905.8]
  wire [57:0] _T_4622; // @[Counters.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@175907.8]
  wire [63:0] _GEN_134; // @[CSR.scala 1058:31:freechips.rocketchip.system.DefaultRV32Config.fir@175903.6]
  wire [31:0] _T_4624; // @[CSR.scala 1059:74:freechips.rocketchip.system.DefaultRV32Config.fir@175912.8]
  wire [63:0] _T_4625; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@175913.8]
  wire [57:0] _T_4626; // @[Counters.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@175915.8]
  wire [63:0] _GEN_136; // @[CSR.scala 1059:31:freechips.rocketchip.system.DefaultRV32Config.fir@175910.6]
  wire [31:0] _T_4627; // @[CSR.scala 1058:47:freechips.rocketchip.system.DefaultRV32Config.fir@175919.8]
  wire [63:0] _T_4628; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@175920.8]
  wire [57:0] _T_4629; // @[Counters.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@175922.8]
  wire [63:0] _GEN_138; // @[CSR.scala 1058:31:freechips.rocketchip.system.DefaultRV32Config.fir@175918.6]
  wire [31:0] _T_4631; // @[CSR.scala 1059:74:freechips.rocketchip.system.DefaultRV32Config.fir@175927.8]
  wire [63:0] _T_4632; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@175928.8]
  wire [57:0] _T_4633; // @[Counters.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@175930.8]
  wire [63:0] _GEN_140; // @[CSR.scala 1059:31:freechips.rocketchip.system.DefaultRV32Config.fir@175925.6]
  wire [31:0] _GEN_143; // @[CSR.scala 858:40:freechips.rocketchip.system.DefaultRV32Config.fir@175933.6]
  wire [31:0] _GEN_145; // @[CSR.scala 859:40:freechips.rocketchip.system.DefaultRV32Config.fir@175937.6]
  wire [26:0] _T_4634; // @[CSR.scala 865:26:freechips.rocketchip.system.DefaultRV32Config.fir@175944.8]
  wire [31:0] _GEN_147; // @[CSR.scala 862:38:freechips.rocketchip.system.DefaultRV32Config.fir@175941.6]
  wire [31:0] _GEN_148; // @[CSR.scala 862:38:freechips.rocketchip.system.DefaultRV32Config.fir@175941.6]
  wire [1:0] _T_4637; // @[CSR.scala 872:43:freechips.rocketchip.system.DefaultRV32Config.fir@175953.8]
  wire  _T_4644; // @[CSR.scala 872:43:freechips.rocketchip.system.DefaultRV32Config.fir@175967.8]
  wire  _T_4647; // @[CSR.scala 872:43:freechips.rocketchip.system.DefaultRV32Config.fir@175973.8]
  wire  _T_4651; // @[CSR.scala 1048:37:freechips.rocketchip.system.DefaultRV32Config.fir@175984.8]
  wire  _T_4658; // @[CSR.scala 924:37:freechips.rocketchip.system.DefaultRV32Config.fir@176005.6]
  wire  _T_4659; // @[CSR.scala 924:55:freechips.rocketchip.system.DefaultRV32Config.fir@176006.6]
  wire  _T_4663; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176018.10]
  wire  _T_4664; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176020.10]
  wire  _T_4666; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176024.10]
  wire  _T_4669; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176030.10]
  wire [1:0] _T_4670; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176032.10]
  wire [31:0] _T_4693; // @[CSR.scala 1043:9:freechips.rocketchip.system.DefaultRV32Config.fir@176064.10]
  wire [31:0] _T_4694; // @[CSR.scala 1043:34:freechips.rocketchip.system.DefaultRV32Config.fir@176065.10]
  wire [31:0] _T_4699; // @[CSR.scala 1043:43:freechips.rocketchip.system.DefaultRV32Config.fir@176070.10]
  wire  _T_4712; // @[CSR.scala 933:96:freechips.rocketchip.system.DefaultRV32Config.fir@176096.10]
  wire  _T_4715; // @[CSR.scala 933:96:freechips.rocketchip.system.DefaultRV32Config.fir@176102.10]
  wire  _T_4717; // @[CSR.scala 934:38:freechips.rocketchip.system.DefaultRV32Config.fir@176106.10]
  wire  _GEN_158; // @[CSR.scala 936:51:freechips.rocketchip.system.DefaultRV32Config.fir@176113.10]
  wire  _T_4801; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176252.6]
  wire  _T_4802; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176253.6]
  wire [7:0] _T_4805; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176258.8 :freechips.rocketchip.system.DefaultRV32Config.fir@176260.8]
  wire  _T_4806; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176261.8]
  wire  _T_4807; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176263.8]
  wire  _T_4808; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176265.8]
  wire [1:0] _T_4809; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176267.8]
  wire  _T_4811; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176271.8]
  wire  _T_4812; // @[CSR.scala 948:31:freechips.rocketchip.system.DefaultRV32Config.fir@176274.8]
  wire  _T_4813; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176277.6]
  wire  _T_4814; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176278.6]
  wire  _T_4816; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176280.6]
  wire  _T_4817; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176281.6]
  wire  _T_4818; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176282.6]
  wire  _T_4819; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176283.6]
  wire  _T_4820; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176284.6]
  wire [31:0] _GEN_229; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176285.6]
  wire  _T_4821; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176288.6]
  wire  _T_4822; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176289.6]
  wire [23:0] _T_4823; // @[CSR.scala 945:53:freechips.rocketchip.system.DefaultRV32Config.fir@176291.8]
  wire [7:0] _T_4825; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176294.8 :freechips.rocketchip.system.DefaultRV32Config.fir@176296.8]
  wire  _T_4826; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176297.8]
  wire  _T_4827; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176299.8]
  wire  _T_4828; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176301.8]
  wire [1:0] _T_4829; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176303.8]
  wire  _T_4831; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176307.8]
  wire  _T_4832; // @[CSR.scala 948:31:freechips.rocketchip.system.DefaultRV32Config.fir@176310.8]
  wire  _T_4833; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176313.6]
  wire  _T_4834; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176314.6]
  wire  _T_4836; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176316.6]
  wire  _T_4837; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176317.6]
  wire  _T_4838; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176318.6]
  wire  _T_4839; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176319.6]
  wire  _T_4840; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176320.6]
  wire [31:0] _GEN_236; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176321.6]
  wire  _T_4841; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176324.6]
  wire  _T_4842; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176325.6]
  wire [15:0] _T_4843; // @[CSR.scala 945:53:freechips.rocketchip.system.DefaultRV32Config.fir@176327.8]
  wire [7:0] _T_4845; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176330.8 :freechips.rocketchip.system.DefaultRV32Config.fir@176332.8]
  wire  _T_4846; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176333.8]
  wire  _T_4847; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176335.8]
  wire  _T_4848; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176337.8]
  wire [1:0] _T_4849; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176339.8]
  wire  _T_4851; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176343.8]
  wire  _T_4852; // @[CSR.scala 948:31:freechips.rocketchip.system.DefaultRV32Config.fir@176346.8]
  wire  _T_4853; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176349.6]
  wire  _T_4854; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176350.6]
  wire  _T_4856; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176352.6]
  wire  _T_4857; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176353.6]
  wire  _T_4858; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176354.6]
  wire  _T_4859; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176355.6]
  wire  _T_4860; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176356.6]
  wire [31:0] _GEN_243; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176357.6]
  wire  _T_4861; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176360.6]
  wire  _T_4862; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176361.6]
  wire [7:0] _T_4863; // @[CSR.scala 945:53:freechips.rocketchip.system.DefaultRV32Config.fir@176363.8]
  wire  _T_4866; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176369.8]
  wire  _T_4867; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176371.8]
  wire  _T_4868; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176373.8]
  wire [1:0] _T_4869; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176375.8]
  wire  _T_4871; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176379.8]
  wire  _T_4872; // @[CSR.scala 948:31:freechips.rocketchip.system.DefaultRV32Config.fir@176382.8]
  wire  _T_4873; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176385.6]
  wire  _T_4874; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176386.6]
  wire  _T_4876; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176388.6]
  wire  _T_4877; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176389.6]
  wire  _T_4878; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176390.6]
  wire  _T_4879; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176391.6]
  wire  _T_4880; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176392.6]
  wire [31:0] _GEN_250; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176393.6]
  wire  _T_4881; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176396.6]
  wire  _T_4882; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176397.6]
  wire  _T_4893; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176421.6]
  wire  _T_4894; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176422.6]
  wire  _T_4896; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176424.6]
  wire  _T_4897; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176425.6]
  wire  _T_4898; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176426.6]
  wire  _T_4899; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176427.6]
  wire  _T_4900; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176428.6]
  wire [31:0] _GEN_257; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176429.6]
  wire  _T_4901; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176432.6]
  wire  _T_4902; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176433.6]
  wire  _T_4913; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176457.6]
  wire  _T_4914; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176458.6]
  wire  _T_4916; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176460.6]
  wire  _T_4917; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176461.6]
  wire  _T_4918; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176462.6]
  wire  _T_4919; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176463.6]
  wire  _T_4920; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176464.6]
  wire [31:0] _GEN_264; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176465.6]
  wire  _T_4921; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176468.6]
  wire  _T_4922; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176469.6]
  wire  _T_4933; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176493.6]
  wire  _T_4934; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176494.6]
  wire  _T_4936; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176496.6]
  wire  _T_4937; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176497.6]
  wire  _T_4938; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176498.6]
  wire  _T_4939; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176499.6]
  wire  _T_4940; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176500.6]
  wire [31:0] _GEN_271; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176501.6]
  wire  _T_4941; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176504.6]
  wire  _T_4942; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176505.6]
  wire  _T_4958; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176534.6]
  wire  _T_4959; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176535.6]
  wire  _T_4960; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176536.6]
  wire [31:0] _GEN_278; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176537.6]
  wire [63:0] _GEN_300; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [63:0] _GEN_302; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_305; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_306; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_353; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_360; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_367; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_374; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_381; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_388; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_395; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire [31:0] _GEN_402; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  wire  _T_5007; // @[CSR.scala 1022:26:freechips.rocketchip.system.DefaultRV32Config.fir@176696.4]
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 574:31:freechips.rocketchip.system.DefaultRV32Config.fir@171058.4]
  assign _T_804 = {io_rw_addr, 20'h0}; // @[CSR.scala 586:28:freechips.rocketchip.system.DefaultRV32Config.fir@171059.4]
  assign _T_811 = _T_804 & 32'h20400000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171066.4]
  assign _T_812 = _T_811 == 32'h20000000; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171067.4]
  assign insn_ret = system_insn & _T_812; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171080.4]
  assign _T_1729 = io_rw_addr[10]; // @[CSR.scala 729:47:freechips.rocketchip.system.DefaultRV32Config.fir@172091.8]
  assign _GEN_93 = _T_1729 ? reg_dcsr_prv : reg_mstatus_mpp; // @[CSR.scala 729:53:freechips.rocketchip.system.DefaultRV32Config.fir@172093.8]
  assign _T_805 = _T_804 & 32'h20100000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171060.4]
  assign _T_806 = _T_805 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171061.4]
  assign insn_call = system_insn & _T_806; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171076.4]
  assign _T_808 = _T_804 & 32'h10100000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171063.4]
  assign _T_809 = _T_808 == 32'h100000; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171064.4]
  assign insn_break = system_insn & _T_809; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171078.4]
  assign _T_1388 = insn_call | insn_break; // @[CSR.scala 658:29:freechips.rocketchip.system.DefaultRV32Config.fir@171680.4]
  assign exception = _T_1388 | io_exception; // @[CSR.scala 658:43:freechips.rocketchip.system.DefaultRV32Config.fir@171681.4]
  assign _GEN_439 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 622:36:freechips.rocketchip.system.DefaultRV32Config.fir@171602.4]
  assign _T_1334 = _GEN_439 + 4'h8; // @[CSR.scala 622:36:freechips.rocketchip.system.DefaultRV32Config.fir@171603.4]
  assign _T_1335 = insn_break ? 32'h3 : io_cause; // @[CSR.scala 623:14:freechips.rocketchip.system.DefaultRV32Config.fir@171604.4]
  assign cause = insn_call ? {{28'd0}, _T_1334} : _T_1335; // @[CSR.scala 622:8:freechips.rocketchip.system.DefaultRV32Config.fir@171605.4]
  assign _T_1336 = cause[31]; // @[CSR.scala 625:30:freechips.rocketchip.system.DefaultRV32Config.fir@171607.4]
  assign cause_lsbs = cause[7:0]; // @[CSR.scala 624:25:freechips.rocketchip.system.DefaultRV32Config.fir@171606.4]
  assign _T_1337 = cause_lsbs == 8'he; // @[CSR.scala 625:53:freechips.rocketchip.system.DefaultRV32Config.fir@171608.4]
  assign causeIsDebugInt = _T_1336 & _T_1337; // @[CSR.scala 625:39:freechips.rocketchip.system.DefaultRV32Config.fir@171609.4]
  assign _T_1349 = reg_singleStepped | causeIsDebugInt; // @[CSR.scala 628:60:freechips.rocketchip.system.DefaultRV32Config.fir@171623.4]
  assign _T_1339 = _T_1336 == 1'h0; // @[CSR.scala 626:29:freechips.rocketchip.system.DefaultRV32Config.fir@171611.4]
  assign causeIsDebugTrigger = _T_1339 & _T_1337; // @[CSR.scala 626:44:freechips.rocketchip.system.DefaultRV32Config.fir@171613.4]
  assign _T_1350 = _T_1349 | causeIsDebugTrigger; // @[CSR.scala 628:79:freechips.rocketchip.system.DefaultRV32Config.fir@171624.4]
  assign _T_1343 = _T_1339 & insn_break; // @[CSR.scala 627:42:freechips.rocketchip.system.DefaultRV32Config.fir@171616.4]
  assign _T_1346 = {reg_dcsr_ebreakm,1'h0,1'h0,reg_dcsr_ebreaku}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@171619.4]
  assign _T_1347 = _T_1346 >> reg_mstatus_prv; // @[CSR.scala 627:134:freechips.rocketchip.system.DefaultRV32Config.fir@171620.4]
  assign _T_1348 = _T_1347[0]; // @[CSR.scala 627:134:freechips.rocketchip.system.DefaultRV32Config.fir@171621.4]
  assign causeIsDebugBreak = _T_1343 & _T_1348; // @[CSR.scala 627:56:freechips.rocketchip.system.DefaultRV32Config.fir@171622.4]
  assign _T_1351 = _T_1350 | causeIsDebugBreak; // @[CSR.scala 628:102:freechips.rocketchip.system.DefaultRV32Config.fir@171625.4]
  assign trapToDebug = _T_1351 | reg_debug; // @[CSR.scala 628:123:freechips.rocketchip.system.DefaultRV32Config.fir@171626.4]
  assign _T_1423 = reg_debug == 1'h0; // @[CSR.scala 675:13:freechips.rocketchip.system.DefaultRV32Config.fir@171746.8]
  assign _GEN_42 = _T_1423 ? 2'h3 : reg_mstatus_prv; // @[CSR.scala 675:25:freechips.rocketchip.system.DefaultRV32Config.fir@171747.8]
  assign _T_1354 = reg_mstatus_prv <= 2'h1; // @[CSR.scala 630:51:freechips.rocketchip.system.DefaultRV32Config.fir@171630.4]
  assign _GEN_61 = trapToDebug ? _GEN_42 : 2'h3; // @[CSR.scala 674:24:freechips.rocketchip.system.DefaultRV32Config.fir@171745.6]
  assign _GEN_79 = exception ? _GEN_61 : reg_mstatus_prv; // @[CSR.scala 673:20:freechips.rocketchip.system.DefaultRV32Config.fir@171744.4]
  assign new_prv = insn_ret ? _GEN_93 : _GEN_79; // @[CSR.scala 722:19:freechips.rocketchip.system.DefaultRV32Config.fir@172074.4]
  assign _T_33 = new_prv[0]; // @[CSR.scala 1048:37:freechips.rocketchip.system.DefaultRV32Config.fir@170129.4]
  assign read_mcounteren = reg_mcounteren & 32'h7; // @[CSR.scala 380:30:freechips.rocketchip.system.DefaultRV32Config.fir@170248.4]
  assign _GEN_440 = {{5'd0}, io_retire}; // @[Counters.scala 47:33:freechips.rocketchip.system.DefaultRV32Config.fir@170263.4]
  assign _T_88 = _T_87 + _GEN_440; // @[Counters.scala 47:33:freechips.rocketchip.system.DefaultRV32Config.fir@170263.4]
  assign _T_90 = _T_88[6]; // @[Counters.scala 52:20:freechips.rocketchip.system.DefaultRV32Config.fir@170266.4]
  assign _T_92 = _T_89 + 58'h1; // @[Counters.scala 52:43:freechips.rocketchip.system.DefaultRV32Config.fir@170269.6]
  assign _T_93 = {_T_89,_T_87}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170272.4]
  assign _T_94 = io_csr_stall == 1'h0; // @[CSR.scala 403:103:freechips.rocketchip.system.DefaultRV32Config.fir@170273.4]
  assign _GEN_441 = {{5'd0}, _T_94}; // @[Counters.scala 47:33:freechips.rocketchip.system.DefaultRV32Config.fir@170275.4]
  assign _T_96 = _T_95 + _GEN_441; // @[Counters.scala 47:33:freechips.rocketchip.system.DefaultRV32Config.fir@170275.4]
  assign _T_98 = _T_96[6]; // @[Counters.scala 52:20:freechips.rocketchip.system.DefaultRV32Config.fir@170278.4]
  assign _T_100 = _T_97 + 58'h1; // @[Counters.scala 52:43:freechips.rocketchip.system.DefaultRV32Config.fir@170281.6]
  assign _T_101 = {_T_97,_T_95}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170284.4]
  assign _T_116 = {4'h0,io_interrupts_meip,1'h0,2'h0,io_interrupts_mtip,1'h0,2'h0,io_interrupts_msip,1'h0,2'h0}; // @[CSR.scala 416:22:freechips.rocketchip.system.DefaultRV32Config.fir@170306.4]
  assign read_mip = _T_116 & 16'h888; // @[CSR.scala 416:29:freechips.rocketchip.system.DefaultRV32Config.fir@170307.4]
  assign _GEN_442 = {{16'd0}, read_mip}; // @[CSR.scala 419:56:freechips.rocketchip.system.DefaultRV32Config.fir@170308.4]
  assign pending_interrupts = _GEN_442 & reg_mie; // @[CSR.scala 419:56:freechips.rocketchip.system.DefaultRV32Config.fir@170308.4]
  assign d_interrupts = {io_interrupts_debug, 14'h0}; // @[CSR.scala 420:42:freechips.rocketchip.system.DefaultRV32Config.fir@170310.4]
  assign _T_119 = _T_1354 | reg_mstatus_mie; // @[CSR.scala 421:51:freechips.rocketchip.system.DefaultRV32Config.fir@170312.4]
  assign _T_120 = ~ pending_interrupts; // @[CSR.scala 421:73:freechips.rocketchip.system.DefaultRV32Config.fir@170313.4]
  assign _T_122 = ~ _T_120; // @[CSR.scala 421:71:freechips.rocketchip.system.DefaultRV32Config.fir@170315.4]
  assign m_interrupts = _T_119 ? _T_122 : 32'h0; // @[CSR.scala 421:25:freechips.rocketchip.system.DefaultRV32Config.fir@170316.4]
  assign _T_128 = d_interrupts[14]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170323.4]
  assign _T_129 = d_interrupts[13]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170324.4]
  assign _T_130 = d_interrupts[12]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170325.4]
  assign _T_131 = d_interrupts[11]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170326.4]
  assign _T_132 = d_interrupts[3]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170327.4]
  assign _T_133 = d_interrupts[7]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170328.4]
  assign _T_134 = d_interrupts[9]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170329.4]
  assign _T_135 = d_interrupts[1]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170330.4]
  assign _T_136 = d_interrupts[5]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170331.4]
  assign _T_137 = d_interrupts[8]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170332.4]
  assign _T_138 = d_interrupts[0]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170333.4]
  assign _T_139 = d_interrupts[4]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170334.4]
  assign _T_140 = m_interrupts[15]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170335.4]
  assign _T_141 = m_interrupts[14]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170336.4]
  assign _T_142 = m_interrupts[13]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170337.4]
  assign _T_143 = m_interrupts[12]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170338.4]
  assign _T_144 = m_interrupts[11]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170339.4]
  assign _T_145 = m_interrupts[3]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170340.4]
  assign _T_146 = m_interrupts[7]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170341.4]
  assign _T_147 = m_interrupts[9]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170342.4]
  assign _T_148 = m_interrupts[1]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170343.4]
  assign _T_149 = m_interrupts[5]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170344.4]
  assign _T_150 = m_interrupts[8]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170345.4]
  assign _T_151 = m_interrupts[0]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170346.4]
  assign _T_152 = m_interrupts[4]; // @[CSR.scala 1037:76:freechips.rocketchip.system.DefaultRV32Config.fir@170347.4]
  assign _T_166 = _T_128 | _T_129; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170361.4]
  assign _T_167 = _T_166 | _T_130; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170362.4]
  assign _T_168 = _T_167 | _T_131; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170363.4]
  assign _T_169 = _T_168 | _T_132; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170364.4]
  assign _T_170 = _T_169 | _T_133; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170365.4]
  assign _T_171 = _T_170 | _T_134; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170366.4]
  assign _T_172 = _T_171 | _T_135; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170367.4]
  assign _T_173 = _T_172 | _T_136; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170368.4]
  assign _T_174 = _T_173 | _T_137; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170369.4]
  assign _T_175 = _T_174 | _T_138; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170370.4]
  assign _T_176 = _T_175 | _T_139; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170371.4]
  assign _T_177 = _T_176 | _T_140; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170372.4]
  assign _T_178 = _T_177 | _T_141; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170373.4]
  assign _T_179 = _T_178 | _T_142; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170374.4]
  assign _T_180 = _T_179 | _T_143; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170375.4]
  assign _T_181 = _T_180 | _T_144; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170376.4]
  assign _T_182 = _T_181 | _T_145; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170377.4]
  assign _T_183 = _T_182 | _T_146; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170378.4]
  assign _T_184 = _T_183 | _T_147; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170379.4]
  assign _T_185 = _T_184 | _T_148; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170380.4]
  assign _T_186 = _T_185 | _T_149; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170381.4]
  assign _T_187 = _T_186 | _T_150; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170382.4]
  assign _T_188 = _T_187 | _T_151; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170383.4]
  assign anyInterrupt = _T_188 | _T_152; // @[CSR.scala 1037:90:freechips.rocketchip.system.DefaultRV32Config.fir@170384.4]
  assign _T_253 = _T_151 ? 4'h0 : 4'h4; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170449.4]
  assign _T_254 = _T_150 ? 4'h8 : _T_253; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170450.4]
  assign _T_255 = _T_149 ? 4'h5 : _T_254; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170451.4]
  assign _T_256 = _T_148 ? 4'h1 : _T_255; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170452.4]
  assign _T_257 = _T_147 ? 4'h9 : _T_256; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170453.4]
  assign _T_258 = _T_146 ? 4'h7 : _T_257; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170454.4]
  assign _T_259 = _T_145 ? 4'h3 : _T_258; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170455.4]
  assign _T_260 = _T_144 ? 4'hb : _T_259; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170456.4]
  assign _T_261 = _T_143 ? 4'hc : _T_260; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170457.4]
  assign _T_262 = _T_142 ? 4'hd : _T_261; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170458.4]
  assign _T_263 = _T_141 ? 4'he : _T_262; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170459.4]
  assign _T_264 = _T_140 ? 4'hf : _T_263; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170460.4]
  assign _T_265 = _T_139 ? 4'h4 : _T_264; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170461.4]
  assign _T_266 = _T_138 ? 4'h0 : _T_265; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170462.4]
  assign _T_267 = _T_137 ? 4'h8 : _T_266; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170463.4]
  assign _T_268 = _T_136 ? 4'h5 : _T_267; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170464.4]
  assign _T_269 = _T_135 ? 4'h1 : _T_268; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170465.4]
  assign _T_270 = _T_134 ? 4'h9 : _T_269; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170466.4]
  assign _T_271 = _T_133 ? 4'h7 : _T_270; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170467.4]
  assign _T_272 = _T_132 ? 4'h3 : _T_271; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170468.4]
  assign _T_273 = _T_131 ? 4'hb : _T_272; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170469.4]
  assign _T_274 = _T_130 ? 4'hc : _T_273; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170470.4]
  assign _T_275 = _T_129 ? 4'hd : _T_274; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170471.4]
  assign whichInterrupt = _T_128 ? 4'he : _T_275; // @[Mux.scala 47:69:freechips.rocketchip.system.DefaultRV32Config.fir@170472.4]
  assign _GEN_443 = {{28'd0}, whichInterrupt}; // @[CSR.scala 425:43:freechips.rocketchip.system.DefaultRV32Config.fir@170473.4]
  assign _T_277 = io_singleStep == 1'h0; // @[CSR.scala 426:36:freechips.rocketchip.system.DefaultRV32Config.fir@170475.4]
  assign _T_278 = anyInterrupt & _T_277; // @[CSR.scala 426:33:freechips.rocketchip.system.DefaultRV32Config.fir@170476.4]
  assign _T_279 = _T_278 | reg_singleStepped; // @[CSR.scala 426:51:freechips.rocketchip.system.DefaultRV32Config.fir@170477.4]
  assign _T_280 = reg_debug | io_status_cease; // @[CSR.scala 426:88:freechips.rocketchip.system.DefaultRV32Config.fir@170478.4]
  assign _T_281 = _T_280 == 1'h0; // @[CSR.scala 426:76:freechips.rocketchip.system.DefaultRV32Config.fir@170479.4]
  assign _T_284 = reg_pmp_0_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170487.4]
  assign _T_285 = {reg_pmp_0_addr,_T_284}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170488.4]
  assign _T_288 = _T_285 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170491.4]
  assign _T_289 = ~ _T_288; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170492.4]
  assign _T_290 = _T_285 & _T_289; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170493.4]
  assign _T_291 = {_T_290,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170494.4]
  assign _T_293 = reg_pmp_1_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170499.4]
  assign _T_294 = {reg_pmp_1_addr,_T_293}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170500.4]
  assign _T_297 = _T_294 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170503.4]
  assign _T_298 = ~ _T_297; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170504.4]
  assign _T_299 = _T_294 & _T_298; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170505.4]
  assign _T_300 = {_T_299,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170506.4]
  assign _T_302 = reg_pmp_2_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170511.4]
  assign _T_303 = {reg_pmp_2_addr,_T_302}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170512.4]
  assign _T_306 = _T_303 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170515.4]
  assign _T_307 = ~ _T_306; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170516.4]
  assign _T_308 = _T_303 & _T_307; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170517.4]
  assign _T_309 = {_T_308,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170518.4]
  assign _T_311 = reg_pmp_3_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170523.4]
  assign _T_312 = {reg_pmp_3_addr,_T_311}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170524.4]
  assign _T_315 = _T_312 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170527.4]
  assign _T_316 = ~ _T_315; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170528.4]
  assign _T_317 = _T_312 & _T_316; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170529.4]
  assign _T_318 = {_T_317,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170530.4]
  assign _T_320 = reg_pmp_4_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170535.4]
  assign _T_321 = {reg_pmp_4_addr,_T_320}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170536.4]
  assign _T_324 = _T_321 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170539.4]
  assign _T_325 = ~ _T_324; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170540.4]
  assign _T_326 = _T_321 & _T_325; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170541.4]
  assign _T_327 = {_T_326,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170542.4]
  assign _T_329 = reg_pmp_5_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170547.4]
  assign _T_330 = {reg_pmp_5_addr,_T_329}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170548.4]
  assign _T_333 = _T_330 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170551.4]
  assign _T_334 = ~ _T_333; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170552.4]
  assign _T_335 = _T_330 & _T_334; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170553.4]
  assign _T_336 = {_T_335,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170554.4]
  assign _T_338 = reg_pmp_6_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170559.4]
  assign _T_339 = {reg_pmp_6_addr,_T_338}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170560.4]
  assign _T_342 = _T_339 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170563.4]
  assign _T_343 = ~ _T_342; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170564.4]
  assign _T_344 = _T_339 & _T_343; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170565.4]
  assign _T_345 = {_T_344,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170566.4]
  assign _T_347 = reg_pmp_7_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.DefaultRV32Config.fir@170571.4]
  assign _T_348 = {reg_pmp_7_addr,_T_347}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170572.4]
  assign _T_351 = _T_348 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.DefaultRV32Config.fir@170575.4]
  assign _T_352 = ~ _T_351; // @[PMP.scala 58:16:freechips.rocketchip.system.DefaultRV32Config.fir@170576.4]
  assign _T_353 = _T_348 & _T_352; // @[PMP.scala 58:14:freechips.rocketchip.system.DefaultRV32Config.fir@170577.4]
  assign _T_354 = {_T_353,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170578.4]
  assign _T_360 = {io_status_hpie,io_status_spie,io_status_upie,io_status_mie,io_status_hie,io_status_sie,io_status_uie}; // @[CSR.scala 445:38:freechips.rocketchip.system.DefaultRV32Config.fir@170594.4]
  assign _T_368 = {io_status_sum,io_status_mprv,io_status_xs,io_status_fs,io_status_mpp,io_status_hpp,io_status_spp,io_status_mpie,_T_360}; // @[CSR.scala 445:38:freechips.rocketchip.system.DefaultRV32Config.fir@170602.4]
  assign _T_375 = {io_status_uxl,io_status_sd_rv32,io_status_zero1,io_status_vs,io_status_tsr,io_status_tw,io_status_tvm,io_status_mxr}; // @[CSR.scala 445:38:freechips.rocketchip.system.DefaultRV32Config.fir@170609.4]
  assign _T_384 = {io_status_debug,io_status_cease,io_status_isa,io_status_dprv,io_status_prv,io_status_sd,io_status_zero2,io_status_sxl,_T_375,_T_368}; // @[CSR.scala 445:38:freechips.rocketchip.system.DefaultRV32Config.fir@170618.4]
  assign read_mstatus = _T_384[31:0]; // @[CSR.scala 445:40:freechips.rocketchip.system.DefaultRV32Config.fir@170619.4]
  assign _T_385 = reg_mtvec[0]; // @[CSR.scala 1066:41:freechips.rocketchip.system.DefaultRV32Config.fir@170620.4]
  assign _T_386 = _T_385 ? 7'h7e : 7'h2; // @[CSR.scala 1066:39:freechips.rocketchip.system.DefaultRV32Config.fir@170621.4]
  assign _T_388 = {{25'd0}, _T_386}; // @[package.scala 131:41:freechips.rocketchip.system.DefaultRV32Config.fir@170623.4]
  assign _T_389 = ~ _T_388; // @[package.scala 131:37:freechips.rocketchip.system.DefaultRV32Config.fir@170624.4]
  assign read_mtvec = reg_mtvec & _T_389; // @[package.scala 131:35:freechips.rocketchip.system.DefaultRV32Config.fir@170625.4]
  assign _T_400 = {reg_bp_0_control_m,1'h0,1'h0,reg_bp_0_control_u,reg_bp_0_control_x,reg_bp_0_control_w,reg_bp_0_control_r}; // @[CSR.scala 451:48:freechips.rocketchip.system.DefaultRV32Config.fir@170637.4]
  assign _T_408 = {4'h2,reg_bp_0_control_dmode,14'h400,reg_bp_0_control_action,1'h0,2'h0,reg_bp_0_control_tmatch,_T_400}; // @[CSR.scala 451:48:freechips.rocketchip.system.DefaultRV32Config.fir@170645.4]
  assign _T_409 = ~ reg_mepc; // @[CSR.scala 1065:28:freechips.rocketchip.system.DefaultRV32Config.fir@170646.4]
  assign _T_410 = reg_misa[2]; // @[CSR.scala 1065:45:freechips.rocketchip.system.DefaultRV32Config.fir@170647.4]
  assign _T_411 = _T_410 ? 2'h1 : 2'h3; // @[CSR.scala 1065:36:freechips.rocketchip.system.DefaultRV32Config.fir@170648.4]
  assign _GEN_444 = {{30'd0}, _T_411}; // @[CSR.scala 1065:31:freechips.rocketchip.system.DefaultRV32Config.fir@170649.4]
  assign _T_412 = _T_409 | _GEN_444; // @[CSR.scala 1065:31:freechips.rocketchip.system.DefaultRV32Config.fir@170649.4]
  assign _T_413 = ~ _T_412; // @[CSR.scala 1065:26:freechips.rocketchip.system.DefaultRV32Config.fir@170650.4]
  assign _T_419 = {2'h0,1'h0,reg_dcsr_cause,3'h0,reg_dcsr_step,reg_dcsr_prv}; // @[CSR.scala 465:27:freechips.rocketchip.system.DefaultRV32Config.fir@170656.4]
  assign _T_426 = {4'h4,12'h0,reg_dcsr_ebreakm,2'h0,reg_dcsr_ebreaku,_T_419}; // @[CSR.scala 465:27:freechips.rocketchip.system.DefaultRV32Config.fir@170663.4]
  assign _T_427 = ~ reg_dpc; // @[CSR.scala 1065:28:freechips.rocketchip.system.DefaultRV32Config.fir@170664.4]
  assign _T_430 = _T_427 | _GEN_444; // @[CSR.scala 1065:31:freechips.rocketchip.system.DefaultRV32Config.fir@170667.4]
  assign _T_431 = ~ _T_430; // @[CSR.scala 1065:26:freechips.rocketchip.system.DefaultRV32Config.fir@170668.4]
  assign _T_432 = {reg_frm,reg_fflags}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170669.4]
  assign _T_434 = {{1'd0}, _T_432}; // @[CSR.scala 469:44:freechips.rocketchip.system.DefaultRV32Config.fir@170671.4]
  assign read_fcsr = {{1'd0}, _T_434}; // @[CSR.scala 469:78:freechips.rocketchip.system.DefaultRV32Config.fir@170673.4]
  assign _T_494 = _T_101[63:32]; // @[CSR.scala 509:50:freechips.rocketchip.system.DefaultRV32Config.fir@170732.4]
  assign _T_495 = _T_93[63:32]; // @[CSR.scala 510:54:freechips.rocketchip.system.DefaultRV32Config.fir@170733.4]
  assign _T_512 = {reg_pmp_0_cfg_l,2'h0,reg_pmp_0_cfg_a,reg_pmp_0_cfg_x,reg_pmp_0_cfg_w,reg_pmp_0_cfg_r}; // @[package.scala 36:38:freechips.rocketchip.system.DefaultRV32Config.fir@170761.4]
  assign _T_522 = {reg_pmp_2_cfg_l,2'h0,reg_pmp_2_cfg_a,reg_pmp_2_cfg_x,reg_pmp_2_cfg_w,reg_pmp_2_cfg_r}; // @[package.scala 36:38:freechips.rocketchip.system.DefaultRV32Config.fir@170771.4]
  assign _T_528 = {reg_pmp_1_cfg_l,2'h0,reg_pmp_1_cfg_a,reg_pmp_1_cfg_x,reg_pmp_1_cfg_w,reg_pmp_1_cfg_r,_T_512}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170777.4]
  assign _T_530 = {reg_pmp_3_cfg_l,2'h0,reg_pmp_3_cfg_a,reg_pmp_3_cfg_x,reg_pmp_3_cfg_w,reg_pmp_3_cfg_r,_T_522,_T_528}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170779.4]
  assign _T_535 = {reg_pmp_4_cfg_l,2'h0,reg_pmp_4_cfg_a,reg_pmp_4_cfg_x,reg_pmp_4_cfg_w,reg_pmp_4_cfg_r}; // @[package.scala 36:38:freechips.rocketchip.system.DefaultRV32Config.fir@170784.4]
  assign _T_545 = {reg_pmp_6_cfg_l,2'h0,reg_pmp_6_cfg_a,reg_pmp_6_cfg_x,reg_pmp_6_cfg_w,reg_pmp_6_cfg_r}; // @[package.scala 36:38:freechips.rocketchip.system.DefaultRV32Config.fir@170794.4]
  assign _T_551 = {reg_pmp_5_cfg_l,2'h0,reg_pmp_5_cfg_a,reg_pmp_5_cfg_x,reg_pmp_5_cfg_w,reg_pmp_5_cfg_r,_T_535}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170800.4]
  assign _T_553 = {reg_pmp_7_cfg_l,2'h0,reg_pmp_7_cfg_a,reg_pmp_7_cfg_x,reg_pmp_7_cfg_w,reg_pmp_7_cfg_r,_T_545,_T_551}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@170802.4]
  assign _T_601 = io_rw_addr == 12'h7a1; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170854.4]
  assign _T_602 = io_rw_addr == 12'h7a2; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170855.4]
  assign _T_603 = io_rw_addr == 12'h301; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170856.4]
  assign _T_604 = io_rw_addr == 12'h300; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170857.4]
  assign _T_605 = io_rw_addr == 12'h305; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170858.4]
  assign _T_606 = io_rw_addr == 12'h344; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170859.4]
  assign _T_607 = io_rw_addr == 12'h304; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170860.4]
  assign _T_608 = io_rw_addr == 12'h340; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170861.4]
  assign _T_609 = io_rw_addr == 12'h341; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170862.4]
  assign _T_610 = io_rw_addr == 12'h343; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170863.4]
  assign _T_611 = io_rw_addr == 12'h342; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170864.4]
  assign _T_613 = io_rw_addr == 12'h7b0; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170866.4]
  assign _T_614 = io_rw_addr == 12'h7b1; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170867.4]
  assign _T_615 = io_rw_addr == 12'h7b2; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170868.4]
  assign _T_616 = io_rw_addr == 12'h1; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170869.4]
  assign _T_617 = io_rw_addr == 12'h2; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170870.4]
  assign _T_618 = io_rw_addr == 12'h3; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170871.4]
  assign _T_619 = io_rw_addr == 12'hb00; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170872.4]
  assign _T_620 = io_rw_addr == 12'hb02; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@170873.4]
  assign _T_766 = io_rw_addr == 12'h306; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171019.4]
  assign _T_767 = io_rw_addr == 12'hc00; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171020.4]
  assign _T_768 = io_rw_addr == 12'hc02; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171021.4]
  assign _T_769 = io_rw_addr == 12'hb80; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171022.4]
  assign _T_770 = io_rw_addr == 12'hb82; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171023.4]
  assign _T_771 = io_rw_addr == 12'hc80; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171024.4]
  assign _T_772 = io_rw_addr == 12'hc82; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171025.4]
  assign _T_773 = io_rw_addr == 12'h3a0; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171026.4]
  assign _T_774 = io_rw_addr == 12'h3a1; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171027.4]
  assign _T_777 = io_rw_addr == 12'h3b0; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171030.4]
  assign _T_778 = io_rw_addr == 12'h3b1; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171031.4]
  assign _T_779 = io_rw_addr == 12'h3b2; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171032.4]
  assign _T_780 = io_rw_addr == 12'h3b3; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171033.4]
  assign _T_781 = io_rw_addr == 12'h3b4; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171034.4]
  assign _T_782 = io_rw_addr == 12'h3b5; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171035.4]
  assign _T_783 = io_rw_addr == 12'h3b6; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171036.4]
  assign _T_784 = io_rw_addr == 12'h3b7; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171037.4]
  assign _T_794 = io_rw_addr == 12'hf12; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171047.4]
  assign _T_796 = io_rw_addr == 12'hf13; // @[CSR.scala 571:73:freechips.rocketchip.system.DefaultRV32Config.fir@171049.4]
  assign _T_797 = io_rw_cmd[1]; // @[CSR.scala 1043:13:freechips.rocketchip.system.DefaultRV32Config.fir@171050.4]
  assign _T_798 = _T_797 ? io_rw_rdata : 32'h0; // @[CSR.scala 1043:9:freechips.rocketchip.system.DefaultRV32Config.fir@171051.4]
  assign _T_799 = _T_798 | io_rw_wdata; // @[CSR.scala 1043:34:freechips.rocketchip.system.DefaultRV32Config.fir@171052.4]
  assign _T_800 = io_rw_cmd[1:0]; // @[CSR.scala 1043:53:freechips.rocketchip.system.DefaultRV32Config.fir@171053.4]
  assign _T_801 = _T_800 == 2'h3; // @[CSR.scala 1043:59:freechips.rocketchip.system.DefaultRV32Config.fir@171054.4]
  assign _T_802 = _T_801 ? io_rw_wdata : 32'h0; // @[CSR.scala 1043:49:freechips.rocketchip.system.DefaultRV32Config.fir@171055.4]
  assign _T_803 = ~ _T_802; // @[CSR.scala 1043:45:freechips.rocketchip.system.DefaultRV32Config.fir@171056.4]
  assign wdata = _T_799 & _T_803; // @[CSR.scala 1043:43:freechips.rocketchip.system.DefaultRV32Config.fir@171057.4]
  assign _T_814 = _T_804 & 32'h20200000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171069.4]
  assign _T_815 = _T_814 == 32'h20000000; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171070.4]
  assign _T_817 = _T_804 & 32'h30000000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171072.4]
  assign _T_818 = _T_817 == 32'h10000000; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171073.4]
  assign insn_cease = system_insn & _T_815; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171082.4]
  assign insn_wfi = system_insn & _T_818; // @[CSR.scala 586:95:freechips.rocketchip.system.DefaultRV32Config.fir@171084.4]
  assign _T_825 = {io_decode_0_csr, 20'h0}; // @[CSR.scala 593:30:freechips.rocketchip.system.DefaultRV32Config.fir@171086.4]
  assign _T_832 = _T_825 & 32'h20400000; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171093.4]
  assign _T_833 = _T_832 == 32'h20000000; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171094.4]
  assign _T_846 = reg_mstatus_prv > 2'h1; // @[CSR.scala 595:55:freechips.rocketchip.system.DefaultRV32Config.fir@171107.4]
  assign _T_858 = io_decode_0_csr[4:0]; // @[CSR.scala 598:34:freechips.rocketchip.system.DefaultRV32Config.fir@171119.4]
  assign _T_860 = read_mcounteren >> _T_858; // @[CSR.scala 599:68:freechips.rocketchip.system.DefaultRV32Config.fir@171121.4]
  assign _T_861 = _T_860[0]; // @[CSR.scala 599:68:freechips.rocketchip.system.DefaultRV32Config.fir@171122.4]
  assign _T_862 = _T_846 | _T_861; // @[CSR.scala 599:50:freechips.rocketchip.system.DefaultRV32Config.fir@171123.4]
  assign _T_869 = io_status_fs == 2'h0; // @[CSR.scala 601:39:freechips.rocketchip.system.DefaultRV32Config.fir@171130.4]
  assign _T_870 = reg_misa[5]; // @[CSR.scala 601:57:freechips.rocketchip.system.DefaultRV32Config.fir@171131.4]
  assign _T_871 = _T_870 == 1'h0; // @[CSR.scala 601:48:freechips.rocketchip.system.DefaultRV32Config.fir@171132.4]
  assign _T_877 = io_decode_0_csr & 12'ha00; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171140.4]
  assign _T_885 = io_decode_0_csr[9:8]; // @[CSR.scala 605:56:freechips.rocketchip.system.DefaultRV32Config.fir@171150.4]
  assign _T_886 = reg_mstatus_prv < _T_885; // @[CSR.scala 605:44:freechips.rocketchip.system.DefaultRV32Config.fir@171151.4]
  assign _T_887 = io_decode_0_csr == 12'h7a0; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171152.4]
  assign _T_888 = io_decode_0_csr == 12'h7a1; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171153.4]
  assign _T_889 = io_decode_0_csr == 12'h7a2; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171154.4]
  assign _T_890 = io_decode_0_csr == 12'h301; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171155.4]
  assign _T_891 = io_decode_0_csr == 12'h300; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171156.4]
  assign _T_892 = io_decode_0_csr == 12'h305; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171157.4]
  assign _T_893 = io_decode_0_csr == 12'h344; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171158.4]
  assign _T_894 = io_decode_0_csr == 12'h304; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171159.4]
  assign _T_895 = io_decode_0_csr == 12'h340; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171160.4]
  assign _T_896 = io_decode_0_csr == 12'h341; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171161.4]
  assign _T_897 = io_decode_0_csr == 12'h343; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171162.4]
  assign _T_898 = io_decode_0_csr == 12'h342; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171163.4]
  assign _T_899 = io_decode_0_csr == 12'hf14; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171164.4]
  assign _T_900 = io_decode_0_csr == 12'h7b0; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171165.4]
  assign _T_901 = io_decode_0_csr == 12'h7b1; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171166.4]
  assign _T_902 = io_decode_0_csr == 12'h7b2; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171167.4]
  assign _T_903 = io_decode_0_csr == 12'h1; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171168.4]
  assign _T_904 = io_decode_0_csr == 12'h2; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171169.4]
  assign _T_905 = io_decode_0_csr == 12'h3; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171170.4]
  assign _T_906 = io_decode_0_csr == 12'hb00; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171171.4]
  assign _T_907 = io_decode_0_csr == 12'hb02; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171172.4]
  assign _T_908 = io_decode_0_csr == 12'h323; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171173.4]
  assign _T_909 = io_decode_0_csr == 12'hb03; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171174.4]
  assign _T_910 = io_decode_0_csr == 12'hc03; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171175.4]
  assign _T_911 = io_decode_0_csr == 12'hb83; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171176.4]
  assign _T_912 = io_decode_0_csr == 12'hc83; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171177.4]
  assign _T_913 = io_decode_0_csr == 12'h324; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171178.4]
  assign _T_914 = io_decode_0_csr == 12'hb04; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171179.4]
  assign _T_915 = io_decode_0_csr == 12'hc04; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171180.4]
  assign _T_916 = io_decode_0_csr == 12'hb84; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171181.4]
  assign _T_917 = io_decode_0_csr == 12'hc84; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171182.4]
  assign _T_918 = io_decode_0_csr == 12'h325; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171183.4]
  assign _T_919 = io_decode_0_csr == 12'hb05; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171184.4]
  assign _T_920 = io_decode_0_csr == 12'hc05; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171185.4]
  assign _T_921 = io_decode_0_csr == 12'hb85; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171186.4]
  assign _T_922 = io_decode_0_csr == 12'hc85; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171187.4]
  assign _T_923 = io_decode_0_csr == 12'h326; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171188.4]
  assign _T_924 = io_decode_0_csr == 12'hb06; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171189.4]
  assign _T_925 = io_decode_0_csr == 12'hc06; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171190.4]
  assign _T_926 = io_decode_0_csr == 12'hb86; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171191.4]
  assign _T_927 = io_decode_0_csr == 12'hc86; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171192.4]
  assign _T_928 = io_decode_0_csr == 12'h327; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171193.4]
  assign _T_929 = io_decode_0_csr == 12'hb07; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171194.4]
  assign _T_930 = io_decode_0_csr == 12'hc07; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171195.4]
  assign _T_931 = io_decode_0_csr == 12'hb87; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171196.4]
  assign _T_932 = io_decode_0_csr == 12'hc87; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171197.4]
  assign _T_933 = io_decode_0_csr == 12'h328; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171198.4]
  assign _T_934 = io_decode_0_csr == 12'hb08; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171199.4]
  assign _T_935 = io_decode_0_csr == 12'hc08; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171200.4]
  assign _T_936 = io_decode_0_csr == 12'hb88; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171201.4]
  assign _T_937 = io_decode_0_csr == 12'hc88; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171202.4]
  assign _T_938 = io_decode_0_csr == 12'h329; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171203.4]
  assign _T_939 = io_decode_0_csr == 12'hb09; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171204.4]
  assign _T_940 = io_decode_0_csr == 12'hc09; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171205.4]
  assign _T_941 = io_decode_0_csr == 12'hb89; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171206.4]
  assign _T_942 = io_decode_0_csr == 12'hc89; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171207.4]
  assign _T_943 = io_decode_0_csr == 12'h32a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171208.4]
  assign _T_944 = io_decode_0_csr == 12'hb0a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171209.4]
  assign _T_945 = io_decode_0_csr == 12'hc0a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171210.4]
  assign _T_946 = io_decode_0_csr == 12'hb8a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171211.4]
  assign _T_947 = io_decode_0_csr == 12'hc8a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171212.4]
  assign _T_948 = io_decode_0_csr == 12'h32b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171213.4]
  assign _T_949 = io_decode_0_csr == 12'hb0b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171214.4]
  assign _T_950 = io_decode_0_csr == 12'hc0b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171215.4]
  assign _T_951 = io_decode_0_csr == 12'hb8b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171216.4]
  assign _T_952 = io_decode_0_csr == 12'hc8b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171217.4]
  assign _T_953 = io_decode_0_csr == 12'h32c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171218.4]
  assign _T_954 = io_decode_0_csr == 12'hb0c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171219.4]
  assign _T_955 = io_decode_0_csr == 12'hc0c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171220.4]
  assign _T_956 = io_decode_0_csr == 12'hb8c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171221.4]
  assign _T_957 = io_decode_0_csr == 12'hc8c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171222.4]
  assign _T_958 = io_decode_0_csr == 12'h32d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171223.4]
  assign _T_959 = io_decode_0_csr == 12'hb0d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171224.4]
  assign _T_960 = io_decode_0_csr == 12'hc0d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171225.4]
  assign _T_961 = io_decode_0_csr == 12'hb8d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171226.4]
  assign _T_962 = io_decode_0_csr == 12'hc8d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171227.4]
  assign _T_963 = io_decode_0_csr == 12'h32e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171228.4]
  assign _T_964 = io_decode_0_csr == 12'hb0e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171229.4]
  assign _T_965 = io_decode_0_csr == 12'hc0e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171230.4]
  assign _T_966 = io_decode_0_csr == 12'hb8e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171231.4]
  assign _T_967 = io_decode_0_csr == 12'hc8e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171232.4]
  assign _T_968 = io_decode_0_csr == 12'h32f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171233.4]
  assign _T_969 = io_decode_0_csr == 12'hb0f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171234.4]
  assign _T_970 = io_decode_0_csr == 12'hc0f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171235.4]
  assign _T_971 = io_decode_0_csr == 12'hb8f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171236.4]
  assign _T_972 = io_decode_0_csr == 12'hc8f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171237.4]
  assign _T_973 = io_decode_0_csr == 12'h330; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171238.4]
  assign _T_974 = io_decode_0_csr == 12'hb10; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171239.4]
  assign _T_975 = io_decode_0_csr == 12'hc10; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171240.4]
  assign _T_976 = io_decode_0_csr == 12'hb90; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171241.4]
  assign _T_977 = io_decode_0_csr == 12'hc90; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171242.4]
  assign _T_978 = io_decode_0_csr == 12'h331; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171243.4]
  assign _T_979 = io_decode_0_csr == 12'hb11; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171244.4]
  assign _T_980 = io_decode_0_csr == 12'hc11; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171245.4]
  assign _T_981 = io_decode_0_csr == 12'hb91; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171246.4]
  assign _T_982 = io_decode_0_csr == 12'hc91; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171247.4]
  assign _T_983 = io_decode_0_csr == 12'h332; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171248.4]
  assign _T_984 = io_decode_0_csr == 12'hb12; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171249.4]
  assign _T_985 = io_decode_0_csr == 12'hc12; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171250.4]
  assign _T_986 = io_decode_0_csr == 12'hb92; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171251.4]
  assign _T_987 = io_decode_0_csr == 12'hc92; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171252.4]
  assign _T_988 = io_decode_0_csr == 12'h333; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171253.4]
  assign _T_989 = io_decode_0_csr == 12'hb13; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171254.4]
  assign _T_990 = io_decode_0_csr == 12'hc13; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171255.4]
  assign _T_991 = io_decode_0_csr == 12'hb93; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171256.4]
  assign _T_992 = io_decode_0_csr == 12'hc93; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171257.4]
  assign _T_993 = io_decode_0_csr == 12'h334; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171258.4]
  assign _T_994 = io_decode_0_csr == 12'hb14; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171259.4]
  assign _T_995 = io_decode_0_csr == 12'hc14; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171260.4]
  assign _T_996 = io_decode_0_csr == 12'hb94; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171261.4]
  assign _T_997 = io_decode_0_csr == 12'hc94; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171262.4]
  assign _T_998 = io_decode_0_csr == 12'h335; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171263.4]
  assign _T_999 = io_decode_0_csr == 12'hb15; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171264.4]
  assign _T_1000 = io_decode_0_csr == 12'hc15; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171265.4]
  assign _T_1001 = io_decode_0_csr == 12'hb95; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171266.4]
  assign _T_1002 = io_decode_0_csr == 12'hc95; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171267.4]
  assign _T_1003 = io_decode_0_csr == 12'h336; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171268.4]
  assign _T_1004 = io_decode_0_csr == 12'hb16; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171269.4]
  assign _T_1005 = io_decode_0_csr == 12'hc16; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171270.4]
  assign _T_1006 = io_decode_0_csr == 12'hb96; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171271.4]
  assign _T_1007 = io_decode_0_csr == 12'hc96; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171272.4]
  assign _T_1008 = io_decode_0_csr == 12'h337; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171273.4]
  assign _T_1009 = io_decode_0_csr == 12'hb17; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171274.4]
  assign _T_1010 = io_decode_0_csr == 12'hc17; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171275.4]
  assign _T_1011 = io_decode_0_csr == 12'hb97; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171276.4]
  assign _T_1012 = io_decode_0_csr == 12'hc97; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171277.4]
  assign _T_1013 = io_decode_0_csr == 12'h338; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171278.4]
  assign _T_1014 = io_decode_0_csr == 12'hb18; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171279.4]
  assign _T_1015 = io_decode_0_csr == 12'hc18; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171280.4]
  assign _T_1016 = io_decode_0_csr == 12'hb98; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171281.4]
  assign _T_1017 = io_decode_0_csr == 12'hc98; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171282.4]
  assign _T_1018 = io_decode_0_csr == 12'h339; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171283.4]
  assign _T_1019 = io_decode_0_csr == 12'hb19; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171284.4]
  assign _T_1020 = io_decode_0_csr == 12'hc19; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171285.4]
  assign _T_1021 = io_decode_0_csr == 12'hb99; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171286.4]
  assign _T_1022 = io_decode_0_csr == 12'hc99; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171287.4]
  assign _T_1023 = io_decode_0_csr == 12'h33a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171288.4]
  assign _T_1024 = io_decode_0_csr == 12'hb1a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171289.4]
  assign _T_1025 = io_decode_0_csr == 12'hc1a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171290.4]
  assign _T_1026 = io_decode_0_csr == 12'hb9a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171291.4]
  assign _T_1027 = io_decode_0_csr == 12'hc9a; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171292.4]
  assign _T_1028 = io_decode_0_csr == 12'h33b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171293.4]
  assign _T_1029 = io_decode_0_csr == 12'hb1b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171294.4]
  assign _T_1030 = io_decode_0_csr == 12'hc1b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171295.4]
  assign _T_1031 = io_decode_0_csr == 12'hb9b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171296.4]
  assign _T_1032 = io_decode_0_csr == 12'hc9b; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171297.4]
  assign _T_1033 = io_decode_0_csr == 12'h33c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171298.4]
  assign _T_1034 = io_decode_0_csr == 12'hb1c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171299.4]
  assign _T_1035 = io_decode_0_csr == 12'hc1c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171300.4]
  assign _T_1036 = io_decode_0_csr == 12'hb9c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171301.4]
  assign _T_1037 = io_decode_0_csr == 12'hc9c; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171302.4]
  assign _T_1038 = io_decode_0_csr == 12'h33d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171303.4]
  assign _T_1039 = io_decode_0_csr == 12'hb1d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171304.4]
  assign _T_1040 = io_decode_0_csr == 12'hc1d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171305.4]
  assign _T_1041 = io_decode_0_csr == 12'hb9d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171306.4]
  assign _T_1042 = io_decode_0_csr == 12'hc9d; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171307.4]
  assign _T_1043 = io_decode_0_csr == 12'h33e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171308.4]
  assign _T_1044 = io_decode_0_csr == 12'hb1e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171309.4]
  assign _T_1045 = io_decode_0_csr == 12'hc1e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171310.4]
  assign _T_1046 = io_decode_0_csr == 12'hb9e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171311.4]
  assign _T_1047 = io_decode_0_csr == 12'hc9e; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171312.4]
  assign _T_1048 = io_decode_0_csr == 12'h33f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171313.4]
  assign _T_1049 = io_decode_0_csr == 12'hb1f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171314.4]
  assign _T_1050 = io_decode_0_csr == 12'hc1f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171315.4]
  assign _T_1051 = io_decode_0_csr == 12'hb9f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171316.4]
  assign _T_1052 = io_decode_0_csr == 12'hc9f; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171317.4]
  assign _T_1053 = io_decode_0_csr == 12'h306; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171318.4]
  assign _T_1054 = io_decode_0_csr == 12'hc00; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171319.4]
  assign _T_1055 = io_decode_0_csr == 12'hc02; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171320.4]
  assign _T_1056 = io_decode_0_csr == 12'hb80; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171321.4]
  assign _T_1057 = io_decode_0_csr == 12'hb82; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171322.4]
  assign _T_1058 = io_decode_0_csr == 12'hc80; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171323.4]
  assign _T_1059 = io_decode_0_csr == 12'hc82; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171324.4]
  assign _T_1060 = io_decode_0_csr == 12'h3a0; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171325.4]
  assign _T_1061 = io_decode_0_csr == 12'h3a1; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171326.4]
  assign _T_1062 = io_decode_0_csr == 12'h3a2; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171327.4]
  assign _T_1063 = io_decode_0_csr == 12'h3a3; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171328.4]
  assign _T_1064 = io_decode_0_csr == 12'h3b0; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171329.4]
  assign _T_1065 = io_decode_0_csr == 12'h3b1; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171330.4]
  assign _T_1066 = io_decode_0_csr == 12'h3b2; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171331.4]
  assign _T_1067 = io_decode_0_csr == 12'h3b3; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171332.4]
  assign _T_1068 = io_decode_0_csr == 12'h3b4; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171333.4]
  assign _T_1069 = io_decode_0_csr == 12'h3b5; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171334.4]
  assign _T_1070 = io_decode_0_csr == 12'h3b6; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171335.4]
  assign _T_1071 = io_decode_0_csr == 12'h3b7; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171336.4]
  assign _T_1072 = io_decode_0_csr == 12'h3b8; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171337.4]
  assign _T_1073 = io_decode_0_csr == 12'h3b9; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171338.4]
  assign _T_1074 = io_decode_0_csr == 12'h3ba; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171339.4]
  assign _T_1075 = io_decode_0_csr == 12'h3bb; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171340.4]
  assign _T_1076 = io_decode_0_csr == 12'h3bc; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171341.4]
  assign _T_1077 = io_decode_0_csr == 12'h3bd; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171342.4]
  assign _T_1078 = io_decode_0_csr == 12'h3be; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171343.4]
  assign _T_1079 = io_decode_0_csr == 12'h3bf; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171344.4]
  assign _T_1080 = io_decode_0_csr == 12'h7c1; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171345.4]
  assign _T_1081 = io_decode_0_csr == 12'hf12; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171346.4]
  assign _T_1082 = io_decode_0_csr == 12'hf11; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171347.4]
  assign _T_1083 = io_decode_0_csr == 12'hf13; // @[CSR.scala 589:99:freechips.rocketchip.system.DefaultRV32Config.fir@171348.4]
  assign _T_1084 = _T_887 | _T_888; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171349.4]
  assign _T_1085 = _T_1084 | _T_889; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171350.4]
  assign _T_1086 = _T_1085 | _T_890; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171351.4]
  assign _T_1087 = _T_1086 | _T_891; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171352.4]
  assign _T_1088 = _T_1087 | _T_892; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171353.4]
  assign _T_1089 = _T_1088 | _T_893; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171354.4]
  assign _T_1090 = _T_1089 | _T_894; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171355.4]
  assign _T_1091 = _T_1090 | _T_895; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171356.4]
  assign _T_1092 = _T_1091 | _T_896; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171357.4]
  assign _T_1093 = _T_1092 | _T_897; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171358.4]
  assign _T_1094 = _T_1093 | _T_898; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171359.4]
  assign _T_1095 = _T_1094 | _T_899; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171360.4]
  assign _T_1096 = _T_1095 | _T_900; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171361.4]
  assign _T_1097 = _T_1096 | _T_901; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171362.4]
  assign _T_1098 = _T_1097 | _T_902; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171363.4]
  assign _T_1099 = _T_1098 | _T_903; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171364.4]
  assign _T_1100 = _T_1099 | _T_904; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171365.4]
  assign _T_1101 = _T_1100 | _T_905; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171366.4]
  assign _T_1102 = _T_1101 | _T_906; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171367.4]
  assign _T_1103 = _T_1102 | _T_907; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171368.4]
  assign _T_1104 = _T_1103 | _T_908; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171369.4]
  assign _T_1105 = _T_1104 | _T_909; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171370.4]
  assign _T_1106 = _T_1105 | _T_910; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171371.4]
  assign _T_1107 = _T_1106 | _T_911; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171372.4]
  assign _T_1108 = _T_1107 | _T_912; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171373.4]
  assign _T_1109 = _T_1108 | _T_913; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171374.4]
  assign _T_1110 = _T_1109 | _T_914; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171375.4]
  assign _T_1111 = _T_1110 | _T_915; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171376.4]
  assign _T_1112 = _T_1111 | _T_916; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171377.4]
  assign _T_1113 = _T_1112 | _T_917; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171378.4]
  assign _T_1114 = _T_1113 | _T_918; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171379.4]
  assign _T_1115 = _T_1114 | _T_919; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171380.4]
  assign _T_1116 = _T_1115 | _T_920; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171381.4]
  assign _T_1117 = _T_1116 | _T_921; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171382.4]
  assign _T_1118 = _T_1117 | _T_922; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171383.4]
  assign _T_1119 = _T_1118 | _T_923; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171384.4]
  assign _T_1120 = _T_1119 | _T_924; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171385.4]
  assign _T_1121 = _T_1120 | _T_925; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171386.4]
  assign _T_1122 = _T_1121 | _T_926; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171387.4]
  assign _T_1123 = _T_1122 | _T_927; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171388.4]
  assign _T_1124 = _T_1123 | _T_928; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171389.4]
  assign _T_1125 = _T_1124 | _T_929; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171390.4]
  assign _T_1126 = _T_1125 | _T_930; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171391.4]
  assign _T_1127 = _T_1126 | _T_931; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171392.4]
  assign _T_1128 = _T_1127 | _T_932; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171393.4]
  assign _T_1129 = _T_1128 | _T_933; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171394.4]
  assign _T_1130 = _T_1129 | _T_934; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171395.4]
  assign _T_1131 = _T_1130 | _T_935; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171396.4]
  assign _T_1132 = _T_1131 | _T_936; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171397.4]
  assign _T_1133 = _T_1132 | _T_937; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171398.4]
  assign _T_1134 = _T_1133 | _T_938; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171399.4]
  assign _T_1135 = _T_1134 | _T_939; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171400.4]
  assign _T_1136 = _T_1135 | _T_940; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171401.4]
  assign _T_1137 = _T_1136 | _T_941; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171402.4]
  assign _T_1138 = _T_1137 | _T_942; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171403.4]
  assign _T_1139 = _T_1138 | _T_943; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171404.4]
  assign _T_1140 = _T_1139 | _T_944; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171405.4]
  assign _T_1141 = _T_1140 | _T_945; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171406.4]
  assign _T_1142 = _T_1141 | _T_946; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171407.4]
  assign _T_1143 = _T_1142 | _T_947; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171408.4]
  assign _T_1144 = _T_1143 | _T_948; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171409.4]
  assign _T_1145 = _T_1144 | _T_949; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171410.4]
  assign _T_1146 = _T_1145 | _T_950; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171411.4]
  assign _T_1147 = _T_1146 | _T_951; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171412.4]
  assign _T_1148 = _T_1147 | _T_952; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171413.4]
  assign _T_1149 = _T_1148 | _T_953; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171414.4]
  assign _T_1150 = _T_1149 | _T_954; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171415.4]
  assign _T_1151 = _T_1150 | _T_955; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171416.4]
  assign _T_1152 = _T_1151 | _T_956; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171417.4]
  assign _T_1153 = _T_1152 | _T_957; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171418.4]
  assign _T_1154 = _T_1153 | _T_958; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171419.4]
  assign _T_1155 = _T_1154 | _T_959; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171420.4]
  assign _T_1156 = _T_1155 | _T_960; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171421.4]
  assign _T_1157 = _T_1156 | _T_961; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171422.4]
  assign _T_1158 = _T_1157 | _T_962; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171423.4]
  assign _T_1159 = _T_1158 | _T_963; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171424.4]
  assign _T_1160 = _T_1159 | _T_964; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171425.4]
  assign _T_1161 = _T_1160 | _T_965; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171426.4]
  assign _T_1162 = _T_1161 | _T_966; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171427.4]
  assign _T_1163 = _T_1162 | _T_967; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171428.4]
  assign _T_1164 = _T_1163 | _T_968; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171429.4]
  assign _T_1165 = _T_1164 | _T_969; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171430.4]
  assign _T_1166 = _T_1165 | _T_970; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171431.4]
  assign _T_1167 = _T_1166 | _T_971; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171432.4]
  assign _T_1168 = _T_1167 | _T_972; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171433.4]
  assign _T_1169 = _T_1168 | _T_973; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171434.4]
  assign _T_1170 = _T_1169 | _T_974; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171435.4]
  assign _T_1171 = _T_1170 | _T_975; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171436.4]
  assign _T_1172 = _T_1171 | _T_976; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171437.4]
  assign _T_1173 = _T_1172 | _T_977; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171438.4]
  assign _T_1174 = _T_1173 | _T_978; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171439.4]
  assign _T_1175 = _T_1174 | _T_979; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171440.4]
  assign _T_1176 = _T_1175 | _T_980; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171441.4]
  assign _T_1177 = _T_1176 | _T_981; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171442.4]
  assign _T_1178 = _T_1177 | _T_982; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171443.4]
  assign _T_1179 = _T_1178 | _T_983; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171444.4]
  assign _T_1180 = _T_1179 | _T_984; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171445.4]
  assign _T_1181 = _T_1180 | _T_985; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171446.4]
  assign _T_1182 = _T_1181 | _T_986; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171447.4]
  assign _T_1183 = _T_1182 | _T_987; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171448.4]
  assign _T_1184 = _T_1183 | _T_988; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171449.4]
  assign _T_1185 = _T_1184 | _T_989; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171450.4]
  assign _T_1186 = _T_1185 | _T_990; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171451.4]
  assign _T_1187 = _T_1186 | _T_991; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171452.4]
  assign _T_1188 = _T_1187 | _T_992; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171453.4]
  assign _T_1189 = _T_1188 | _T_993; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171454.4]
  assign _T_1190 = _T_1189 | _T_994; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171455.4]
  assign _T_1191 = _T_1190 | _T_995; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171456.4]
  assign _T_1192 = _T_1191 | _T_996; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171457.4]
  assign _T_1193 = _T_1192 | _T_997; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171458.4]
  assign _T_1194 = _T_1193 | _T_998; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171459.4]
  assign _T_1195 = _T_1194 | _T_999; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171460.4]
  assign _T_1196 = _T_1195 | _T_1000; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171461.4]
  assign _T_1197 = _T_1196 | _T_1001; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171462.4]
  assign _T_1198 = _T_1197 | _T_1002; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171463.4]
  assign _T_1199 = _T_1198 | _T_1003; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171464.4]
  assign _T_1200 = _T_1199 | _T_1004; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171465.4]
  assign _T_1201 = _T_1200 | _T_1005; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171466.4]
  assign _T_1202 = _T_1201 | _T_1006; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171467.4]
  assign _T_1203 = _T_1202 | _T_1007; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171468.4]
  assign _T_1204 = _T_1203 | _T_1008; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171469.4]
  assign _T_1205 = _T_1204 | _T_1009; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171470.4]
  assign _T_1206 = _T_1205 | _T_1010; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171471.4]
  assign _T_1207 = _T_1206 | _T_1011; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171472.4]
  assign _T_1208 = _T_1207 | _T_1012; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171473.4]
  assign _T_1209 = _T_1208 | _T_1013; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171474.4]
  assign _T_1210 = _T_1209 | _T_1014; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171475.4]
  assign _T_1211 = _T_1210 | _T_1015; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171476.4]
  assign _T_1212 = _T_1211 | _T_1016; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171477.4]
  assign _T_1213 = _T_1212 | _T_1017; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171478.4]
  assign _T_1214 = _T_1213 | _T_1018; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171479.4]
  assign _T_1215 = _T_1214 | _T_1019; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171480.4]
  assign _T_1216 = _T_1215 | _T_1020; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171481.4]
  assign _T_1217 = _T_1216 | _T_1021; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171482.4]
  assign _T_1218 = _T_1217 | _T_1022; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171483.4]
  assign _T_1219 = _T_1218 | _T_1023; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171484.4]
  assign _T_1220 = _T_1219 | _T_1024; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171485.4]
  assign _T_1221 = _T_1220 | _T_1025; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171486.4]
  assign _T_1222 = _T_1221 | _T_1026; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171487.4]
  assign _T_1223 = _T_1222 | _T_1027; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171488.4]
  assign _T_1224 = _T_1223 | _T_1028; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171489.4]
  assign _T_1225 = _T_1224 | _T_1029; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171490.4]
  assign _T_1226 = _T_1225 | _T_1030; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171491.4]
  assign _T_1227 = _T_1226 | _T_1031; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171492.4]
  assign _T_1228 = _T_1227 | _T_1032; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171493.4]
  assign _T_1229 = _T_1228 | _T_1033; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171494.4]
  assign _T_1230 = _T_1229 | _T_1034; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171495.4]
  assign _T_1231 = _T_1230 | _T_1035; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171496.4]
  assign _T_1232 = _T_1231 | _T_1036; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171497.4]
  assign _T_1233 = _T_1232 | _T_1037; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171498.4]
  assign _T_1234 = _T_1233 | _T_1038; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171499.4]
  assign _T_1235 = _T_1234 | _T_1039; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171500.4]
  assign _T_1236 = _T_1235 | _T_1040; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171501.4]
  assign _T_1237 = _T_1236 | _T_1041; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171502.4]
  assign _T_1238 = _T_1237 | _T_1042; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171503.4]
  assign _T_1239 = _T_1238 | _T_1043; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171504.4]
  assign _T_1240 = _T_1239 | _T_1044; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171505.4]
  assign _T_1241 = _T_1240 | _T_1045; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171506.4]
  assign _T_1242 = _T_1241 | _T_1046; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171507.4]
  assign _T_1243 = _T_1242 | _T_1047; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171508.4]
  assign _T_1244 = _T_1243 | _T_1048; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171509.4]
  assign _T_1245 = _T_1244 | _T_1049; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171510.4]
  assign _T_1246 = _T_1245 | _T_1050; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171511.4]
  assign _T_1247 = _T_1246 | _T_1051; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171512.4]
  assign _T_1248 = _T_1247 | _T_1052; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171513.4]
  assign _T_1249 = _T_1248 | _T_1053; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171514.4]
  assign _T_1250 = _T_1249 | _T_1054; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171515.4]
  assign _T_1251 = _T_1250 | _T_1055; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171516.4]
  assign _T_1252 = _T_1251 | _T_1056; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171517.4]
  assign _T_1253 = _T_1252 | _T_1057; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171518.4]
  assign _T_1254 = _T_1253 | _T_1058; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171519.4]
  assign _T_1255 = _T_1254 | _T_1059; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171520.4]
  assign _T_1256 = _T_1255 | _T_1060; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171521.4]
  assign _T_1257 = _T_1256 | _T_1061; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171522.4]
  assign _T_1258 = _T_1257 | _T_1062; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171523.4]
  assign _T_1259 = _T_1258 | _T_1063; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171524.4]
  assign _T_1260 = _T_1259 | _T_1064; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171525.4]
  assign _T_1261 = _T_1260 | _T_1065; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171526.4]
  assign _T_1262 = _T_1261 | _T_1066; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171527.4]
  assign _T_1263 = _T_1262 | _T_1067; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171528.4]
  assign _T_1264 = _T_1263 | _T_1068; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171529.4]
  assign _T_1265 = _T_1264 | _T_1069; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171530.4]
  assign _T_1266 = _T_1265 | _T_1070; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171531.4]
  assign _T_1267 = _T_1266 | _T_1071; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171532.4]
  assign _T_1268 = _T_1267 | _T_1072; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171533.4]
  assign _T_1269 = _T_1268 | _T_1073; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171534.4]
  assign _T_1270 = _T_1269 | _T_1074; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171535.4]
  assign _T_1271 = _T_1270 | _T_1075; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171536.4]
  assign _T_1272 = _T_1271 | _T_1076; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171537.4]
  assign _T_1273 = _T_1272 | _T_1077; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171538.4]
  assign _T_1274 = _T_1273 | _T_1078; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171539.4]
  assign _T_1275 = _T_1274 | _T_1079; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171540.4]
  assign _T_1276 = _T_1275 | _T_1080; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171541.4]
  assign _T_1277 = _T_1276 | _T_1081; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171542.4]
  assign _T_1278 = _T_1277 | _T_1082; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171543.4]
  assign _T_1279 = _T_1278 | _T_1083; // @[CSR.scala 589:115:freechips.rocketchip.system.DefaultRV32Config.fir@171544.4]
  assign _T_1280 = _T_1279 == 1'h0; // @[CSR.scala 606:7:freechips.rocketchip.system.DefaultRV32Config.fir@171545.4]
  assign _T_1281 = _T_886 | _T_1280; // @[CSR.scala 605:62:freechips.rocketchip.system.DefaultRV32Config.fir@171546.4]
  assign _T_1286 = io_decode_0_csr >= 12'hc00; // @[package.scala 162:47:freechips.rocketchip.system.DefaultRV32Config.fir@171551.4]
  assign _T_1287 = io_decode_0_csr < 12'hc20; // @[package.scala 162:60:freechips.rocketchip.system.DefaultRV32Config.fir@171552.4]
  assign _T_1288 = _T_1286 & _T_1287; // @[package.scala 162:55:freechips.rocketchip.system.DefaultRV32Config.fir@171553.4]
  assign _T_1289 = io_decode_0_csr >= 12'hc80; // @[package.scala 162:47:freechips.rocketchip.system.DefaultRV32Config.fir@171554.4]
  assign _T_1290 = io_decode_0_csr < 12'hca0; // @[package.scala 162:60:freechips.rocketchip.system.DefaultRV32Config.fir@171555.4]
  assign _T_1291 = _T_1289 & _T_1290; // @[package.scala 162:55:freechips.rocketchip.system.DefaultRV32Config.fir@171556.4]
  assign _T_1292 = _T_1288 | _T_1291; // @[CSR.scala 608:66:freechips.rocketchip.system.DefaultRV32Config.fir@171557.4]
  assign _T_1293 = _T_862 == 1'h0; // @[CSR.scala 608:133:freechips.rocketchip.system.DefaultRV32Config.fir@171558.4]
  assign _T_1294 = _T_1292 & _T_1293; // @[CSR.scala 608:130:freechips.rocketchip.system.DefaultRV32Config.fir@171559.4]
  assign _T_1295 = _T_1281 | _T_1294; // @[CSR.scala 607:53:freechips.rocketchip.system.DefaultRV32Config.fir@171560.4]
  assign _T_1296 = io_decode_0_csr & 12'hc10; // @[Decode.scala 14:65:freechips.rocketchip.system.DefaultRV32Config.fir@171561.4]
  assign _T_1297 = _T_1296 == 12'h410; // @[Decode.scala 14:121:freechips.rocketchip.system.DefaultRV32Config.fir@171562.4]
  assign _T_1301 = _T_1297 & _T_1423; // @[CSR.scala 609:42:freechips.rocketchip.system.DefaultRV32Config.fir@171566.4]
  assign _T_1302 = _T_1295 | _T_1301; // @[CSR.scala 608:148:freechips.rocketchip.system.DefaultRV32Config.fir@171567.4]
  assign _T_1305 = io_decode_0_fp_csr & io_decode_0_fp_illegal; // @[CSR.scala 611:21:freechips.rocketchip.system.DefaultRV32Config.fir@171570.4]
  assign _T_1307 = io_decode_0_csr[11:10]; // @[CSR.scala 612:39:freechips.rocketchip.system.DefaultRV32Config.fir@171573.4]
  assign _T_1309 = io_decode_0_csr >= 12'h340; // @[CSR.scala 613:40:freechips.rocketchip.system.DefaultRV32Config.fir@171576.4]
  assign _T_1310 = io_decode_0_csr <= 12'h343; // @[CSR.scala 613:71:freechips.rocketchip.system.DefaultRV32Config.fir@171577.4]
  assign _T_1311 = _T_1309 & _T_1310; // @[CSR.scala 613:57:freechips.rocketchip.system.DefaultRV32Config.fir@171578.4]
  assign _T_1312 = io_decode_0_csr >= 12'h140; // @[CSR.scala 613:99:freechips.rocketchip.system.DefaultRV32Config.fir@171579.4]
  assign _T_1313 = io_decode_0_csr <= 12'h143; // @[CSR.scala 613:130:freechips.rocketchip.system.DefaultRV32Config.fir@171580.4]
  assign _T_1314 = _T_1312 & _T_1313; // @[CSR.scala 613:116:freechips.rocketchip.system.DefaultRV32Config.fir@171581.4]
  assign _T_1315 = _T_1311 | _T_1314; // @[CSR.scala 613:85:freechips.rocketchip.system.DefaultRV32Config.fir@171582.4]
  assign _T_1325 = io_decode_0_csr[10]; // @[CSR.scala 617:27:freechips.rocketchip.system.DefaultRV32Config.fir@171593.4]
  assign _T_1326 = _T_833 & _T_1325; // @[CSR.scala 617:14:freechips.rocketchip.system.DefaultRV32Config.fir@171594.4]
  assign _T_1328 = _T_1326 & _T_1423; // @[CSR.scala 617:32:freechips.rocketchip.system.DefaultRV32Config.fir@171596.4]
  assign _T_1353 = insn_break ? 12'h800 : 12'h808; // @[CSR.scala 629:37:freechips.rocketchip.system.DefaultRV32Config.fir@171628.4]
  assign debugTVec = reg_debug ? _T_1353 : 12'h800; // @[CSR.scala 629:22:freechips.rocketchip.system.DefaultRV32Config.fir@171629.4]
  assign _T_1363 = cause[4:0]; // @[CSR.scala 638:32:freechips.rocketchip.system.DefaultRV32Config.fir@171640.4]
  assign _T_1364 = {_T_1363, 2'h0}; // @[CSR.scala 638:59:freechips.rocketchip.system.DefaultRV32Config.fir@171641.4]
  assign _T_1365 = read_mtvec[31:7]; // @[CSR.scala 639:33:freechips.rocketchip.system.DefaultRV32Config.fir@171642.4]
  assign _T_1366 = {_T_1365,_T_1364}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@171643.4]
  assign _T_1367 = read_mtvec[0]; // @[CSR.scala 640:24:freechips.rocketchip.system.DefaultRV32Config.fir@171644.4]
  assign _T_1369 = _T_1367 & _T_1336; // @[CSR.scala 640:28:freechips.rocketchip.system.DefaultRV32Config.fir@171646.4]
  assign _T_1370 = cause_lsbs[7:5]; // @[CSR.scala 640:70:freechips.rocketchip.system.DefaultRV32Config.fir@171647.4]
  assign _T_1371 = _T_1370 == 3'h0; // @[CSR.scala 640:94:freechips.rocketchip.system.DefaultRV32Config.fir@171648.4]
  assign _T_1372 = _T_1369 & _T_1371; // @[CSR.scala 640:55:freechips.rocketchip.system.DefaultRV32Config.fir@171649.4]
  assign _T_1373 = read_mtvec[31:2]; // @[CSR.scala 641:38:freechips.rocketchip.system.DefaultRV32Config.fir@171650.4]
  assign _T_1374 = {_T_1373, 2'h0}; // @[CSR.scala 641:56:freechips.rocketchip.system.DefaultRV32Config.fir@171651.4]
  assign notDebugTVec = _T_1372 ? _T_1366 : _T_1374; // @[CSR.scala 641:8:freechips.rocketchip.system.DefaultRV32Config.fir@171652.4]
  assign tvec = trapToDebug ? {{20'd0}, debugTVec} : notDebugTVec; // @[CSR.scala 643:17:freechips.rocketchip.system.DefaultRV32Config.fir@171653.4]
  assign _T_1379 = io_status_fs == 2'h3; // @[CSR.scala 649:32:freechips.rocketchip.system.DefaultRV32Config.fir@171663.4]
  assign _T_1380 = io_status_xs == 2'h3; // @[CSR.scala 649:53:freechips.rocketchip.system.DefaultRV32Config.fir@171664.4]
  assign _T_1381 = _T_1379 | _T_1380; // @[CSR.scala 649:37:freechips.rocketchip.system.DefaultRV32Config.fir@171665.4]
  assign _T_1382 = io_status_vs == 2'h3; // @[CSR.scala 649:74:freechips.rocketchip.system.DefaultRV32Config.fir@171666.4]
  assign _T_1385 = reg_mstatus_mprv & _T_1423; // @[CSR.scala 654:53:freechips.rocketchip.system.DefaultRV32Config.fir@171674.4]
  assign _T_1389 = insn_ret + insn_call; // @[Bitwise.scala 47:55:freechips.rocketchip.system.DefaultRV32Config.fir@171682.4]
  assign _T_1391 = insn_break + io_exception; // @[Bitwise.scala 47:55:freechips.rocketchip.system.DefaultRV32Config.fir@171684.4]
  assign _T_1393 = _T_1389 + _T_1391; // @[Bitwise.scala 47:55:freechips.rocketchip.system.DefaultRV32Config.fir@171686.4]
  assign _T_1395 = _T_1393 <= 3'h1; // @[CSR.scala 659:79:freechips.rocketchip.system.DefaultRV32Config.fir@171688.4]
  assign _T_1397 = _T_1395 | reset; // @[CSR.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@171690.4]
  assign _T_1398 = _T_1397 == 1'h0; // @[CSR.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@171691.4]
  assign _T_1400 = insn_wfi & _T_277; // @[CSR.scala 661:18:freechips.rocketchip.system.DefaultRV32Config.fir@171697.4]
  assign _T_1402 = _T_1400 & _T_1423; // @[CSR.scala 661:36:freechips.rocketchip.system.DefaultRV32Config.fir@171699.4]
  assign _GEN_34 = _T_1402 | reg_wfi; // @[CSR.scala 661:51:freechips.rocketchip.system.DefaultRV32Config.fir@171700.4]
  assign _T_1403 = pending_interrupts != 32'h0; // @[CSR.scala 662:28:freechips.rocketchip.system.DefaultRV32Config.fir@171703.4]
  assign _T_1404 = _T_1403 | io_interrupts_debug; // @[CSR.scala 662:32:freechips.rocketchip.system.DefaultRV32Config.fir@171704.4]
  assign _T_1405 = _T_1404 | exception; // @[CSR.scala 662:55:freechips.rocketchip.system.DefaultRV32Config.fir@171705.4]
  assign _T_1407 = io_retire | exception; // @[CSR.scala 664:22:freechips.rocketchip.system.DefaultRV32Config.fir@171710.4]
  assign _GEN_36 = _T_1407 | reg_singleStepped; // @[CSR.scala 664:36:freechips.rocketchip.system.DefaultRV32Config.fir@171711.4]
  assign _T_1415 = reg_singleStepped == 1'h0; // @[CSR.scala 667:10:freechips.rocketchip.system.DefaultRV32Config.fir@171728.4]
  assign _T_1416 = io_retire == 1'h0; // @[CSR.scala 667:42:freechips.rocketchip.system.DefaultRV32Config.fir@171729.4]
  assign _T_1417 = _T_1415 | _T_1416; // @[CSR.scala 667:29:freechips.rocketchip.system.DefaultRV32Config.fir@171730.4]
  assign _T_1419 = _T_1417 | reset; // @[CSR.scala 667:9:freechips.rocketchip.system.DefaultRV32Config.fir@171732.4]
  assign _T_1420 = _T_1419 == 1'h0; // @[CSR.scala 667:9:freechips.rocketchip.system.DefaultRV32Config.fir@171733.4]
  assign _T_1421 = ~ io_pc; // @[CSR.scala 1064:28:freechips.rocketchip.system.DefaultRV32Config.fir@171738.4]
  assign _T_1422 = _T_1421 | 32'h1; // @[CSR.scala 1064:31:freechips.rocketchip.system.DefaultRV32Config.fir@171739.4]
  assign epc = ~ _T_1422; // @[CSR.scala 1064:26:freechips.rocketchip.system.DefaultRV32Config.fir@171740.4]
  assign _T_1424 = causeIsDebugTrigger ? 2'h2 : 2'h1; // @[CSR.scala 678:86:freechips.rocketchip.system.DefaultRV32Config.fir@171750.10]
  assign _T_1425 = causeIsDebugInt ? 2'h3 : _T_1424; // @[CSR.scala 678:56:freechips.rocketchip.system.DefaultRV32Config.fir@171751.10]
  assign _T_1427 = reg_mstatus_prv[0]; // @[CSR.scala 1048:37:freechips.rocketchip.system.DefaultRV32Config.fir@171754.10]
  assign _T_1429 = _T_1427 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@171756.10]
  assign _GEN_38 = _T_1423 | reg_debug; // @[CSR.scala 675:25:freechips.rocketchip.system.DefaultRV32Config.fir@171747.8]
  assign _GEN_48 = {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 682:27:freechips.rocketchip.system.DefaultRV32Config.fir@171762.8]
  assign _GEN_67 = trapToDebug ? {{1'd0}, reg_mstatus_spp} : _GEN_48; // @[CSR.scala 674:24:freechips.rocketchip.system.DefaultRV32Config.fir@171745.6]
  assign _GEN_74 = trapToDebug & reg_mstatus_mie; // @[CSR.scala 674:24:freechips.rocketchip.system.DefaultRV32Config.fir@171745.6]
  assign _GEN_85 = exception ? _GEN_67 : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 673:20:freechips.rocketchip.system.DefaultRV32Config.fir@171744.4]
  assign _GEN_95 = _T_1729 ? _T_431 : _T_413; // @[CSR.scala 729:53:freechips.rocketchip.system.DefaultRV32Config.fir@172093.8]
  assign _GEN_117 = insn_cease | _T_1743; // @[Reg.scala 28:19:freechips.rocketchip.system.DefaultRV32Config.fir@172121.4]
  assign _T_1745 = _T_601 ? _T_408 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172138.4]
  assign _T_1746 = _T_602 ? reg_bp_0_address : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172139.4]
  assign _T_1747 = _T_603 ? reg_misa : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172140.4]
  assign _T_1748 = _T_604 ? read_mstatus : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172141.4]
  assign _T_1749 = _T_605 ? read_mtvec : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172142.4]
  assign _T_1750 = _T_606 ? read_mip : 16'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172143.4]
  assign _T_1751 = _T_607 ? reg_mie : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172144.4]
  assign _T_1752 = _T_608 ? reg_mscratch : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172145.4]
  assign _T_1753 = _T_609 ? _T_413 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172146.4]
  assign _T_1754 = _T_610 ? reg_mtval : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172147.4]
  assign _T_1755 = _T_611 ? reg_mcause : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172148.4]
  assign _T_1757 = _T_613 ? _T_426 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172150.4]
  assign _T_1758 = _T_614 ? _T_431 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172151.4]
  assign _T_1759 = _T_615 ? reg_dscratch : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172152.4]
  assign _T_1760 = _T_616 ? reg_fflags : 5'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172153.4]
  assign _T_1761 = _T_617 ? reg_frm : 3'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172154.4]
  assign _T_1762 = _T_618 ? read_fcsr : 10'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172155.4]
  assign _T_1763 = _T_619 ? _T_101 : 64'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172156.4]
  assign _T_1764 = _T_620 ? _T_93 : 64'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172157.4]
  assign _T_1910 = _T_766 ? read_mcounteren : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172303.4]
  assign _T_1911 = _T_767 ? _T_101 : 64'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172304.4]
  assign _T_1912 = _T_768 ? _T_93 : 64'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172305.4]
  assign _T_1913 = _T_769 ? _T_494 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172306.4]
  assign _T_1914 = _T_770 ? _T_495 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172307.4]
  assign _T_1915 = _T_771 ? _T_494 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172308.4]
  assign _T_1916 = _T_772 ? _T_495 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172309.4]
  assign _T_1917 = _T_773 ? _T_530 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172310.4]
  assign _T_1918 = _T_774 ? _T_553 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172311.4]
  assign _T_1921 = _T_777 ? reg_pmp_0_addr : 30'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172314.4]
  assign _T_1922 = _T_778 ? reg_pmp_1_addr : 30'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172315.4]
  assign _T_1923 = _T_779 ? reg_pmp_2_addr : 30'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172316.4]
  assign _T_1924 = _T_780 ? reg_pmp_3_addr : 30'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172317.4]
  assign _T_1925 = _T_781 ? reg_pmp_4_addr : 30'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172318.4]
  assign _T_1926 = _T_782 ? reg_pmp_5_addr : 30'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172319.4]
  assign _T_1927 = _T_783 ? reg_pmp_6_addr : 30'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172320.4]
  assign _T_1928 = _T_784 ? reg_pmp_7_addr : 30'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172321.4]
  assign _T_1938 = _T_794 ? 32'h1 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172331.4]
  assign _T_1940 = _T_796 ? 32'h20181004 : 32'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172333.4]
  assign _T_1942 = _T_1745 | _T_1746; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172335.4]
  assign _T_1943 = _T_1942 | _T_1747; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172336.4]
  assign _T_1944 = _T_1943 | _T_1748; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172337.4]
  assign _T_1945 = _T_1944 | _T_1749; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172338.4]
  assign _GEN_448 = {{16'd0}, _T_1750}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172339.4]
  assign _T_1946 = _T_1945 | _GEN_448; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172339.4]
  assign _T_1947 = _T_1946 | _T_1751; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172340.4]
  assign _T_1948 = _T_1947 | _T_1752; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172341.4]
  assign _T_1949 = _T_1948 | _T_1753; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172342.4]
  assign _T_1950 = _T_1949 | _T_1754; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172343.4]
  assign _T_1951 = _T_1950 | _T_1755; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172344.4]
  assign _T_1953 = _T_1951 | _T_1757; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172346.4]
  assign _T_1954 = _T_1953 | _T_1758; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172347.4]
  assign _T_1955 = _T_1954 | _T_1759; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172348.4]
  assign _GEN_449 = {{27'd0}, _T_1760}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172349.4]
  assign _T_1956 = _T_1955 | _GEN_449; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172349.4]
  assign _GEN_450 = {{29'd0}, _T_1761}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172350.4]
  assign _T_1957 = _T_1956 | _GEN_450; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172350.4]
  assign _GEN_451 = {{22'd0}, _T_1762}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172351.4]
  assign _T_1958 = _T_1957 | _GEN_451; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172351.4]
  assign _GEN_452 = {{32'd0}, _T_1958}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172352.4]
  assign _T_1959 = _GEN_452 | _T_1763; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172352.4]
  assign _T_1960 = _T_1959 | _T_1764; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172353.4]
  assign _GEN_453 = {{32'd0}, _T_1910}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172499.4]
  assign _T_2106 = _T_1960 | _GEN_453; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172499.4]
  assign _T_2107 = _T_2106 | _T_1911; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172500.4]
  assign _T_2108 = _T_2107 | _T_1912; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172501.4]
  assign _GEN_454 = {{32'd0}, _T_1913}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172502.4]
  assign _T_2109 = _T_2108 | _GEN_454; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172502.4]
  assign _GEN_455 = {{32'd0}, _T_1914}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172503.4]
  assign _T_2110 = _T_2109 | _GEN_455; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172503.4]
  assign _GEN_456 = {{32'd0}, _T_1915}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172504.4]
  assign _T_2111 = _T_2110 | _GEN_456; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172504.4]
  assign _GEN_457 = {{32'd0}, _T_1916}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172505.4]
  assign _T_2112 = _T_2111 | _GEN_457; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172505.4]
  assign _GEN_458 = {{32'd0}, _T_1917}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172506.4]
  assign _T_2113 = _T_2112 | _GEN_458; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172506.4]
  assign _GEN_459 = {{32'd0}, _T_1918}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172507.4]
  assign _T_2114 = _T_2113 | _GEN_459; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172507.4]
  assign _GEN_460 = {{34'd0}, _T_1921}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172510.4]
  assign _T_2117 = _T_2114 | _GEN_460; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172510.4]
  assign _GEN_461 = {{34'd0}, _T_1922}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172511.4]
  assign _T_2118 = _T_2117 | _GEN_461; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172511.4]
  assign _GEN_462 = {{34'd0}, _T_1923}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172512.4]
  assign _T_2119 = _T_2118 | _GEN_462; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172512.4]
  assign _GEN_463 = {{34'd0}, _T_1924}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172513.4]
  assign _T_2120 = _T_2119 | _GEN_463; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172513.4]
  assign _GEN_464 = {{34'd0}, _T_1925}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172514.4]
  assign _T_2121 = _T_2120 | _GEN_464; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172514.4]
  assign _GEN_465 = {{34'd0}, _T_1926}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172515.4]
  assign _T_2122 = _T_2121 | _GEN_465; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172515.4]
  assign _GEN_466 = {{34'd0}, _T_1927}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172516.4]
  assign _T_2123 = _T_2122 | _GEN_466; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172516.4]
  assign _GEN_467 = {{34'd0}, _T_1928}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172517.4]
  assign _T_2124 = _T_2123 | _GEN_467; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172517.4]
  assign _GEN_468 = {{32'd0}, _T_1938}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172527.4]
  assign _T_2134 = _T_2124 | _GEN_468; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172527.4]
  assign _GEN_469 = {{32'd0}, _T_1940}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172529.4]
  assign _T_2136 = _T_2134 | _GEN_469; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@172529.4]
  assign _T_2140 = io_rw_cmd == 3'h5; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@172536.6]
  assign _T_2141 = io_rw_cmd == 3'h6; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@172537.6]
  assign _T_2142 = io_rw_cmd == 3'h7; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@172538.6]
  assign _T_4502 = reg_fflags | io_fcsr_flags_bits; // @[CSR.scala 781:30:freechips.rocketchip.system.DefaultRV32Config.fir@175693.6]
  assign _GEN_118 = io_fcsr_flags_valid ? _T_4502 : reg_fflags; // @[CSR.scala 780:30:freechips.rocketchip.system.DefaultRV32Config.fir@175692.4]
  assign _T_4506 = _T_2141 | _T_2142; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@175700.4]
  assign csr_wen = _T_4506 | _T_2140; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@175701.4]
  assign _T_4520 = {{70'd0}, wdata}; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@175719.8 :freechips.rocketchip.system.DefaultRV32Config.fir@175721.8]
  assign _T_4524 = _T_4520[3]; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175728.8]
  assign _T_4528 = _T_4520[7]; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175736.8]
  assign _T_4531 = _T_4520[12:11]; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175742.8]
  assign _T_4532 = _T_4520[14:13]; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175744.8]
  assign _T_4534 = _T_4520[17]; // @[CSR.scala 796:47:freechips.rocketchip.system.DefaultRV32Config.fir@175748.8]
  assign _T_4552 = _T_4531[0]; // @[CSR.scala 1048:37:freechips.rocketchip.system.DefaultRV32Config.fir@175787.8]
  assign _T_4555 = _T_4532 != 2'h0; // @[CSR.scala 1068:73:freechips.rocketchip.system.DefaultRV32Config.fir@175791.8]
  assign _T_4558 = wdata[5]; // @[CSR.scala 821:20:freechips.rocketchip.system.DefaultRV32Config.fir@175798.8]
  assign _T_4559 = io_pc[1]; // @[CSR.scala 823:39:freechips.rocketchip.system.DefaultRV32Config.fir@175799.8]
  assign _T_4560 = _T_4559 == 1'h0; // @[CSR.scala 823:33:freechips.rocketchip.system.DefaultRV32Config.fir@175800.8]
  assign _T_4562 = wdata[2]; // @[CSR.scala 823:51:freechips.rocketchip.system.DefaultRV32Config.fir@175802.8]
  assign _T_4563 = _T_4560 | _T_4562; // @[CSR.scala 823:43:freechips.rocketchip.system.DefaultRV32Config.fir@175803.8]
  assign _T_4564 = ~ wdata; // @[CSR.scala 825:25:freechips.rocketchip.system.DefaultRV32Config.fir@175805.10]
  assign _T_4565 = _T_4558 == 1'h0; // @[CSR.scala 825:35:freechips.rocketchip.system.DefaultRV32Config.fir@175806.10]
  assign _T_4566 = {_T_4565, 3'h0}; // @[CSR.scala 825:38:freechips.rocketchip.system.DefaultRV32Config.fir@175807.10]
  assign _GEN_470 = {{28'd0}, _T_4566}; // @[CSR.scala 825:32:freechips.rocketchip.system.DefaultRV32Config.fir@175808.10]
  assign _T_4567 = _T_4564 | _GEN_470; // @[CSR.scala 825:32:freechips.rocketchip.system.DefaultRV32Config.fir@175808.10]
  assign _T_4568 = ~ _T_4567; // @[CSR.scala 825:23:freechips.rocketchip.system.DefaultRV32Config.fir@175809.10]
  assign _T_4569 = _T_4568 & 32'h1025; // @[CSR.scala 825:55:freechips.rocketchip.system.DefaultRV32Config.fir@175810.10]
  assign _T_4571 = reg_misa & 32'hffffefda; // @[CSR.scala 825:73:freechips.rocketchip.system.DefaultRV32Config.fir@175812.10]
  assign _T_4572 = _T_4569 | _T_4571; // @[CSR.scala 825:62:freechips.rocketchip.system.DefaultRV32Config.fir@175813.10]
  assign _T_4614 = wdata & 32'h888; // @[CSR.scala 840:59:freechips.rocketchip.system.DefaultRV32Config.fir@175880.8]
  assign _T_4616 = _T_4564 | 32'h1; // @[CSR.scala 1064:31:freechips.rocketchip.system.DefaultRV32Config.fir@175885.8]
  assign _T_4617 = ~ _T_4616; // @[CSR.scala 1064:26:freechips.rocketchip.system.DefaultRV32Config.fir@175886.8]
  assign _T_4618 = wdata & 32'h8000000f; // @[CSR.scala 845:62:freechips.rocketchip.system.DefaultRV32Config.fir@175896.8]
  assign _T_4620 = _T_101[63:32]; // @[CSR.scala 1058:47:freechips.rocketchip.system.DefaultRV32Config.fir@175904.8]
  assign _T_4621 = {_T_4620,wdata}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@175905.8]
  assign _T_4622 = _T_4621[63:6]; // @[Counters.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@175907.8]
  assign _GEN_134 = _T_619 ? _T_4621 : {{57'd0}, _T_96}; // @[CSR.scala 1058:31:freechips.rocketchip.system.DefaultRV32Config.fir@175903.6]
  assign _T_4624 = _T_101[31:0]; // @[CSR.scala 1059:74:freechips.rocketchip.system.DefaultRV32Config.fir@175912.8]
  assign _T_4625 = {wdata,_T_4624}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@175913.8]
  assign _T_4626 = _T_4625[63:6]; // @[Counters.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@175915.8]
  assign _GEN_136 = _T_769 ? _T_4625 : _GEN_134; // @[CSR.scala 1059:31:freechips.rocketchip.system.DefaultRV32Config.fir@175910.6]
  assign _T_4627 = _T_93[63:32]; // @[CSR.scala 1058:47:freechips.rocketchip.system.DefaultRV32Config.fir@175919.8]
  assign _T_4628 = {_T_4627,wdata}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@175920.8]
  assign _T_4629 = _T_4628[63:6]; // @[Counters.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@175922.8]
  assign _GEN_138 = _T_620 ? _T_4628 : {{57'd0}, _T_88}; // @[CSR.scala 1058:31:freechips.rocketchip.system.DefaultRV32Config.fir@175918.6]
  assign _T_4631 = _T_93[31:0]; // @[CSR.scala 1059:74:freechips.rocketchip.system.DefaultRV32Config.fir@175927.8]
  assign _T_4632 = {wdata,_T_4631}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@175928.8]
  assign _T_4633 = _T_4632[63:6]; // @[Counters.scala 67:28:freechips.rocketchip.system.DefaultRV32Config.fir@175930.8]
  assign _GEN_140 = _T_770 ? _T_4632 : _GEN_138; // @[CSR.scala 1059:31:freechips.rocketchip.system.DefaultRV32Config.fir@175925.6]
  assign _GEN_143 = _T_616 ? wdata : {{27'd0}, _GEN_118}; // @[CSR.scala 858:40:freechips.rocketchip.system.DefaultRV32Config.fir@175933.6]
  assign _GEN_145 = _T_617 ? wdata : {{29'd0}, reg_frm}; // @[CSR.scala 859:40:freechips.rocketchip.system.DefaultRV32Config.fir@175937.6]
  assign _T_4634 = wdata[31:5]; // @[CSR.scala 865:26:freechips.rocketchip.system.DefaultRV32Config.fir@175944.8]
  assign _GEN_147 = _T_618 ? wdata : _GEN_143; // @[CSR.scala 862:38:freechips.rocketchip.system.DefaultRV32Config.fir@175941.6]
  assign _GEN_148 = _T_618 ? {{5'd0}, _T_4634} : _GEN_145; // @[CSR.scala 862:38:freechips.rocketchip.system.DefaultRV32Config.fir@175941.6]
  assign _T_4637 = wdata[1:0]; // @[CSR.scala 872:43:freechips.rocketchip.system.DefaultRV32Config.fir@175953.8]
  assign _T_4644 = wdata[12]; // @[CSR.scala 872:43:freechips.rocketchip.system.DefaultRV32Config.fir@175967.8]
  assign _T_4647 = wdata[15]; // @[CSR.scala 872:43:freechips.rocketchip.system.DefaultRV32Config.fir@175973.8]
  assign _T_4651 = _T_4637[0]; // @[CSR.scala 1048:37:freechips.rocketchip.system.DefaultRV32Config.fir@175984.8]
  assign _T_4658 = reg_bp_0_control_dmode == 1'h0; // @[CSR.scala 924:37:freechips.rocketchip.system.DefaultRV32Config.fir@176005.6]
  assign _T_4659 = _T_4658 | reg_debug; // @[CSR.scala 924:55:freechips.rocketchip.system.DefaultRV32Config.fir@176006.6]
  assign _T_4663 = wdata[0]; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176018.10]
  assign _T_4664 = wdata[1]; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176020.10]
  assign _T_4666 = wdata[3]; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176024.10]
  assign _T_4669 = wdata[6]; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176030.10]
  assign _T_4670 = wdata[8:7]; // @[CSR.scala 927:41:freechips.rocketchip.system.DefaultRV32Config.fir@176032.10]
  assign _T_4693 = _T_797 ? _T_408 : 32'h0; // @[CSR.scala 1043:9:freechips.rocketchip.system.DefaultRV32Config.fir@176064.10]
  assign _T_4694 = _T_4693 | io_rw_wdata; // @[CSR.scala 1043:34:freechips.rocketchip.system.DefaultRV32Config.fir@176065.10]
  assign _T_4699 = _T_4694 & _T_803; // @[CSR.scala 1043:43:freechips.rocketchip.system.DefaultRV32Config.fir@176070.10]
  assign _T_4712 = _T_4699[12]; // @[CSR.scala 933:96:freechips.rocketchip.system.DefaultRV32Config.fir@176096.10]
  assign _T_4715 = _T_4699[27]; // @[CSR.scala 933:96:freechips.rocketchip.system.DefaultRV32Config.fir@176102.10]
  assign _T_4717 = _T_4715 & reg_debug; // @[CSR.scala 934:38:freechips.rocketchip.system.DefaultRV32Config.fir@176106.10]
  assign _GEN_158 = _T_4717 & _T_4712; // @[CSR.scala 936:51:freechips.rocketchip.system.DefaultRV32Config.fir@176113.10]
  assign _T_4801 = reg_pmp_0_cfg_l == 1'h0; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176252.6]
  assign _T_4802 = _T_773 & _T_4801; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176253.6]
  assign _T_4805 = wdata[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176258.8 :freechips.rocketchip.system.DefaultRV32Config.fir@176260.8]
  assign _T_4806 = _T_4805[0]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176261.8]
  assign _T_4807 = _T_4805[1]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176263.8]
  assign _T_4808 = _T_4805[2]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176265.8]
  assign _T_4809 = _T_4805[4:3]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176267.8]
  assign _T_4811 = _T_4805[7]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176271.8]
  assign _T_4812 = _T_4807 & _T_4806; // @[CSR.scala 948:31:freechips.rocketchip.system.DefaultRV32Config.fir@176274.8]
  assign _T_4813 = reg_pmp_1_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176277.6]
  assign _T_4814 = _T_4813 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176278.6]
  assign _T_4816 = _T_4814 & _T_293; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176280.6]
  assign _T_4817 = reg_pmp_1_cfg_l & _T_4816; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176281.6]
  assign _T_4818 = reg_pmp_0_cfg_l | _T_4817; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176282.6]
  assign _T_4819 = _T_4818 == 1'h0; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176283.6]
  assign _T_4820 = _T_777 & _T_4819; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176284.6]
  assign _GEN_229 = _T_4820 ? wdata : {{2'd0}, reg_pmp_0_addr}; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176285.6]
  assign _T_4821 = reg_pmp_1_cfg_l == 1'h0; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176288.6]
  assign _T_4822 = _T_773 & _T_4821; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176289.6]
  assign _T_4823 = wdata[31:8]; // @[CSR.scala 945:53:freechips.rocketchip.system.DefaultRV32Config.fir@176291.8]
  assign _T_4825 = _T_4823[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176294.8 :freechips.rocketchip.system.DefaultRV32Config.fir@176296.8]
  assign _T_4826 = _T_4825[0]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176297.8]
  assign _T_4827 = _T_4825[1]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176299.8]
  assign _T_4828 = _T_4825[2]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176301.8]
  assign _T_4829 = _T_4825[4:3]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176303.8]
  assign _T_4831 = _T_4825[7]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176307.8]
  assign _T_4832 = _T_4827 & _T_4826; // @[CSR.scala 948:31:freechips.rocketchip.system.DefaultRV32Config.fir@176310.8]
  assign _T_4833 = reg_pmp_2_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176313.6]
  assign _T_4834 = _T_4833 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176314.6]
  assign _T_4836 = _T_4834 & _T_302; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176316.6]
  assign _T_4837 = reg_pmp_2_cfg_l & _T_4836; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176317.6]
  assign _T_4838 = reg_pmp_1_cfg_l | _T_4837; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176318.6]
  assign _T_4839 = _T_4838 == 1'h0; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176319.6]
  assign _T_4840 = _T_778 & _T_4839; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176320.6]
  assign _GEN_236 = _T_4840 ? wdata : {{2'd0}, reg_pmp_1_addr}; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176321.6]
  assign _T_4841 = reg_pmp_2_cfg_l == 1'h0; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176324.6]
  assign _T_4842 = _T_773 & _T_4841; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176325.6]
  assign _T_4843 = wdata[31:16]; // @[CSR.scala 945:53:freechips.rocketchip.system.DefaultRV32Config.fir@176327.8]
  assign _T_4845 = _T_4843[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@176330.8 :freechips.rocketchip.system.DefaultRV32Config.fir@176332.8]
  assign _T_4846 = _T_4845[0]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176333.8]
  assign _T_4847 = _T_4845[1]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176335.8]
  assign _T_4848 = _T_4845[2]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176337.8]
  assign _T_4849 = _T_4845[4:3]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176339.8]
  assign _T_4851 = _T_4845[7]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176343.8]
  assign _T_4852 = _T_4847 & _T_4846; // @[CSR.scala 948:31:freechips.rocketchip.system.DefaultRV32Config.fir@176346.8]
  assign _T_4853 = reg_pmp_3_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176349.6]
  assign _T_4854 = _T_4853 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176350.6]
  assign _T_4856 = _T_4854 & _T_311; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176352.6]
  assign _T_4857 = reg_pmp_3_cfg_l & _T_4856; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176353.6]
  assign _T_4858 = reg_pmp_2_cfg_l | _T_4857; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176354.6]
  assign _T_4859 = _T_4858 == 1'h0; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176355.6]
  assign _T_4860 = _T_779 & _T_4859; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176356.6]
  assign _GEN_243 = _T_4860 ? wdata : {{2'd0}, reg_pmp_2_addr}; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176357.6]
  assign _T_4861 = reg_pmp_3_cfg_l == 1'h0; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176360.6]
  assign _T_4862 = _T_773 & _T_4861; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176361.6]
  assign _T_4863 = wdata[31:24]; // @[CSR.scala 945:53:freechips.rocketchip.system.DefaultRV32Config.fir@176363.8]
  assign _T_4866 = _T_4863[0]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176369.8]
  assign _T_4867 = _T_4863[1]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176371.8]
  assign _T_4868 = _T_4863[2]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176373.8]
  assign _T_4869 = _T_4863[4:3]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176375.8]
  assign _T_4871 = _T_4863[7]; // @[CSR.scala 945:46:freechips.rocketchip.system.DefaultRV32Config.fir@176379.8]
  assign _T_4872 = _T_4867 & _T_4866; // @[CSR.scala 948:31:freechips.rocketchip.system.DefaultRV32Config.fir@176382.8]
  assign _T_4873 = reg_pmp_4_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176385.6]
  assign _T_4874 = _T_4873 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176386.6]
  assign _T_4876 = _T_4874 & _T_320; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176388.6]
  assign _T_4877 = reg_pmp_4_cfg_l & _T_4876; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176389.6]
  assign _T_4878 = reg_pmp_3_cfg_l | _T_4877; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176390.6]
  assign _T_4879 = _T_4878 == 1'h0; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176391.6]
  assign _T_4880 = _T_780 & _T_4879; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176392.6]
  assign _GEN_250 = _T_4880 ? wdata : {{2'd0}, reg_pmp_3_addr}; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176393.6]
  assign _T_4881 = reg_pmp_4_cfg_l == 1'h0; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176396.6]
  assign _T_4882 = _T_774 & _T_4881; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176397.6]
  assign _T_4893 = reg_pmp_5_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176421.6]
  assign _T_4894 = _T_4893 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176422.6]
  assign _T_4896 = _T_4894 & _T_329; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176424.6]
  assign _T_4897 = reg_pmp_5_cfg_l & _T_4896; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176425.6]
  assign _T_4898 = reg_pmp_4_cfg_l | _T_4897; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176426.6]
  assign _T_4899 = _T_4898 == 1'h0; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176427.6]
  assign _T_4900 = _T_781 & _T_4899; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176428.6]
  assign _GEN_257 = _T_4900 ? wdata : {{2'd0}, reg_pmp_4_addr}; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176429.6]
  assign _T_4901 = reg_pmp_5_cfg_l == 1'h0; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176432.6]
  assign _T_4902 = _T_774 & _T_4901; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176433.6]
  assign _T_4913 = reg_pmp_6_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176457.6]
  assign _T_4914 = _T_4913 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176458.6]
  assign _T_4916 = _T_4914 & _T_338; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176460.6]
  assign _T_4917 = reg_pmp_6_cfg_l & _T_4916; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176461.6]
  assign _T_4918 = reg_pmp_5_cfg_l | _T_4917; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176462.6]
  assign _T_4919 = _T_4918 == 1'h0; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176463.6]
  assign _T_4920 = _T_782 & _T_4919; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176464.6]
  assign _GEN_264 = _T_4920 ? wdata : {{2'd0}, reg_pmp_5_addr}; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176465.6]
  assign _T_4921 = reg_pmp_6_cfg_l == 1'h0; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176468.6]
  assign _T_4922 = _T_774 & _T_4921; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176469.6]
  assign _T_4933 = reg_pmp_7_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@176493.6]
  assign _T_4934 = _T_4933 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.DefaultRV32Config.fir@176494.6]
  assign _T_4936 = _T_4934 & _T_347; // @[PMP.scala 47:20:freechips.rocketchip.system.DefaultRV32Config.fir@176496.6]
  assign _T_4937 = reg_pmp_7_cfg_l & _T_4936; // @[PMP.scala 49:62:freechips.rocketchip.system.DefaultRV32Config.fir@176497.6]
  assign _T_4938 = reg_pmp_6_cfg_l | _T_4937; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176498.6]
  assign _T_4939 = _T_4938 == 1'h0; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176499.6]
  assign _T_4940 = _T_783 & _T_4939; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176500.6]
  assign _GEN_271 = _T_4940 ? wdata : {{2'd0}, reg_pmp_6_addr}; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176501.6]
  assign _T_4941 = reg_pmp_7_cfg_l == 1'h0; // @[CSR.scala 944:60:freechips.rocketchip.system.DefaultRV32Config.fir@176504.6]
  assign _T_4942 = _T_774 & _T_4941; // @[CSR.scala 944:57:freechips.rocketchip.system.DefaultRV32Config.fir@176505.6]
  assign _T_4958 = reg_pmp_7_cfg_l | _T_4937; // @[PMP.scala 49:44:freechips.rocketchip.system.DefaultRV32Config.fir@176534.6]
  assign _T_4959 = _T_4958 == 1'h0; // @[CSR.scala 953:48:freechips.rocketchip.system.DefaultRV32Config.fir@176535.6]
  assign _T_4960 = _T_784 & _T_4959; // @[CSR.scala 953:45:freechips.rocketchip.system.DefaultRV32Config.fir@176536.6]
  assign _GEN_278 = _T_4960 ? wdata : {{2'd0}, reg_pmp_7_addr}; // @[CSR.scala 953:71:freechips.rocketchip.system.DefaultRV32Config.fir@176537.6]
  assign _GEN_300 = csr_wen ? _GEN_136 : {{57'd0}, _T_96}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_302 = csr_wen ? _GEN_140 : {{57'd0}, _T_88}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_305 = csr_wen ? _GEN_147 : {{27'd0}, _GEN_118}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_306 = csr_wen ? _GEN_148 : {{29'd0}, reg_frm}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_353 = csr_wen ? _GEN_229 : {{2'd0}, reg_pmp_0_addr}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_360 = csr_wen ? _GEN_236 : {{2'd0}, reg_pmp_1_addr}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_367 = csr_wen ? _GEN_243 : {{2'd0}, reg_pmp_2_addr}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_374 = csr_wen ? _GEN_250 : {{2'd0}, reg_pmp_3_addr}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_381 = csr_wen ? _GEN_257 : {{2'd0}, reg_pmp_4_addr}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_388 = csr_wen ? _GEN_264 : {{2'd0}, reg_pmp_5_addr}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_395 = csr_wen ? _GEN_271 : {{2'd0}, reg_pmp_6_addr}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _GEN_402 = csr_wen ? _GEN_278 : {{2'd0}, reg_pmp_7_addr}; // @[CSR.scala 794:18:freechips.rocketchip.system.DefaultRV32Config.fir@175715.4]
  assign _T_5007 = io_retire > 1'h0; // @[CSR.scala 1022:26:freechips.rocketchip.system.DefaultRV32Config.fir@176696.4]
  assign io_rw_rdata = _T_2136[31:0]; // @[CSR.scala 752:15:freechips.rocketchip.system.DefaultRV32Config.fir@172532.4]
  assign io_decode_0_fp_illegal = _T_869 | _T_871; // @[CSR.scala 601:23:freechips.rocketchip.system.DefaultRV32Config.fir@171134.4]
  assign io_decode_0_fp_csr = _T_877 == 12'h0; // @[CSR.scala 603:19:freechips.rocketchip.system.DefaultRV32Config.fir@171144.4]
  assign io_decode_0_read_illegal = _T_1302 | _T_1305; // @[CSR.scala 605:25:freechips.rocketchip.system.DefaultRV32Config.fir@171572.4]
  assign io_decode_0_write_illegal = _T_1307 == 2'h3; // @[CSR.scala 612:26:freechips.rocketchip.system.DefaultRV32Config.fir@171575.4]
  assign io_decode_0_write_flush = _T_1315 == 1'h0; // @[CSR.scala 613:24:freechips.rocketchip.system.DefaultRV32Config.fir@171584.4]
  assign io_decode_0_system_illegal = _T_886 | _T_1328; // @[CSR.scala 614:27:freechips.rocketchip.system.DefaultRV32Config.fir@171601.4]
  assign io_csr_stall = reg_wfi | io_status_cease; // @[CSR.scala 743:16:freechips.rocketchip.system.DefaultRV32Config.fir@172119.4]
  assign io_eret = _T_1388 | insn_ret; // @[CSR.scala 646:11:freechips.rocketchip.system.DefaultRV32Config.fir@171658.4]
  assign io_singleStep = reg_dcsr_step & _T_1423; // @[CSR.scala 647:17:freechips.rocketchip.system.DefaultRV32Config.fir@171661.4]
  assign io_status_debug = reg_debug; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4 CSR.scala 650:19:freechips.rocketchip.system.DefaultRV32Config.fir@171669.4]
  assign io_status_cease = _T_1743; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4 CSR.scala 744:19:freechips.rocketchip.system.DefaultRV32Config.fir@172124.4]
  assign io_status_isa = reg_misa; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4 CSR.scala 651:17:freechips.rocketchip.system.DefaultRV32Config.fir@171670.4]
  assign io_status_dprv = _T_1387; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4 CSR.scala 654:18:freechips.rocketchip.system.DefaultRV32Config.fir@171678.4]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_sd = _T_1381 | _T_1382; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4 CSR.scala 649:16:freechips.rocketchip.system.DefaultRV32Config.fir@171668.4]
  assign io_status_zero2 = 27'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_sxl = 2'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4 CSR.scala 653:17:freechips.rocketchip.system.DefaultRV32Config.fir@171672.4]
  assign io_status_uxl = 2'h1; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4 CSR.scala 652:17:freechips.rocketchip.system.DefaultRV32Config.fir@171671.4]
  assign io_status_sd_rv32 = io_status_sd; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4 CSR.scala 656:23:freechips.rocketchip.system.DefaultRV32Config.fir@171679.4]
  assign io_status_zero1 = 6'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_vs = 2'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_tsr = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_tw = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_tvm = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_mxr = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_sum = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_mprv = reg_mstatus_mprv; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_xs = 2'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_fs = reg_mstatus_fs; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_mpp = reg_mstatus_mpp; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_hpp = 2'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_spp = reg_mstatus_spp; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_hpie = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_spie = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_upie = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_hie = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_sie = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_status_uie = 1'h0; // @[CSR.scala 648:13:freechips.rocketchip.system.DefaultRV32Config.fir@171662.4]
  assign io_evec = insn_ret ? _GEN_95 : tvec; // @[CSR.scala 644:11:freechips.rocketchip.system.DefaultRV32Config.fir@171654.4 CSR.scala 728:15:freechips.rocketchip.system.DefaultRV32Config.fir@172088.8 CSR.scala 732:15:freechips.rocketchip.system.DefaultRV32Config.fir@172101.10 CSR.scala 738:15:freechips.rocketchip.system.DefaultRV32Config.fir@172114.10]
  assign io_time = _T_101[31:0]; // @[CSR.scala 742:11:freechips.rocketchip.system.DefaultRV32Config.fir@172117.4]
  assign io_fcsr_rm = reg_frm; // @[CSR.scala 779:14:freechips.rocketchip.system.DefaultRV32Config.fir@175691.4]
  assign io_interrupt = _T_279 & _T_281; // @[CSR.scala 426:16:freechips.rocketchip.system.DefaultRV32Config.fir@170481.4]
  assign io_interrupt_cause = 32'h80000000 + _GEN_443; // @[CSR.scala 427:22:freechips.rocketchip.system.DefaultRV32Config.fir@170482.4]
  assign io_bp_0_control_action = reg_bp_0_control_action; // @[CSR.scala 428:9:freechips.rocketchip.system.DefaultRV32Config.fir@170483.4]
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch; // @[CSR.scala 428:9:freechips.rocketchip.system.DefaultRV32Config.fir@170483.4]
  assign io_bp_0_control_m = reg_bp_0_control_m; // @[CSR.scala 428:9:freechips.rocketchip.system.DefaultRV32Config.fir@170483.4]
  assign io_bp_0_control_u = reg_bp_0_control_u; // @[CSR.scala 428:9:freechips.rocketchip.system.DefaultRV32Config.fir@170483.4]
  assign io_bp_0_control_x = reg_bp_0_control_x; // @[CSR.scala 428:9:freechips.rocketchip.system.DefaultRV32Config.fir@170483.4]
  assign io_bp_0_control_w = reg_bp_0_control_w; // @[CSR.scala 428:9:freechips.rocketchip.system.DefaultRV32Config.fir@170483.4]
  assign io_bp_0_control_r = reg_bp_0_control_r; // @[CSR.scala 428:9:freechips.rocketchip.system.DefaultRV32Config.fir@170483.4]
  assign io_bp_0_address = reg_bp_0_address; // @[CSR.scala 428:9:freechips.rocketchip.system.DefaultRV32Config.fir@170483.4]
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170580.4]
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170580.4]
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170580.4]
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170580.4]
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170580.4]
  assign io_pmp_0_addr = reg_pmp_0_addr; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170580.4]
  assign io_pmp_0_mask = _T_291[31:0]; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170580.4]
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170581.4]
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170581.4]
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170581.4]
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170581.4]
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170581.4]
  assign io_pmp_1_addr = reg_pmp_1_addr; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170581.4]
  assign io_pmp_1_mask = _T_300[31:0]; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170581.4]
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170582.4]
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170582.4]
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170582.4]
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170582.4]
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170582.4]
  assign io_pmp_2_addr = reg_pmp_2_addr; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170582.4]
  assign io_pmp_2_mask = _T_309[31:0]; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170582.4]
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170583.4]
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170583.4]
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170583.4]
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170583.4]
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170583.4]
  assign io_pmp_3_addr = reg_pmp_3_addr; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170583.4]
  assign io_pmp_3_mask = _T_318[31:0]; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170583.4]
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170584.4]
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170584.4]
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170584.4]
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170584.4]
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170584.4]
  assign io_pmp_4_addr = reg_pmp_4_addr; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170584.4]
  assign io_pmp_4_mask = _T_327[31:0]; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170584.4]
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170585.4]
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170585.4]
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170585.4]
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170585.4]
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170585.4]
  assign io_pmp_5_addr = reg_pmp_5_addr; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170585.4]
  assign io_pmp_5_mask = _T_336[31:0]; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170585.4]
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170586.4]
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170586.4]
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170586.4]
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170586.4]
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170586.4]
  assign io_pmp_6_addr = reg_pmp_6_addr; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170586.4]
  assign io_pmp_6_mask = _T_345[31:0]; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170586.4]
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170587.4]
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170587.4]
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170587.4]
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170587.4]
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170587.4]
  assign io_pmp_7_addr = reg_pmp_7_addr; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170587.4]
  assign io_pmp_7_mask = _T_354[31:0]; // @[CSR.scala 429:10:freechips.rocketchip.system.DefaultRV32Config.fir@170587.4]
  assign io_trace_0_valid = _T_5007 | io_trace_0_exception; // @[CSR.scala 1022:13:freechips.rocketchip.system.DefaultRV32Config.fir@176698.4]
  assign io_trace_0_iaddr = io_pc; // @[CSR.scala 1024:13:freechips.rocketchip.system.DefaultRV32Config.fir@176700.4]
  assign io_trace_0_insn = io_inst_0; // @[CSR.scala 1023:12:freechips.rocketchip.system.DefaultRV32Config.fir@176699.4]
  assign io_trace_0_exception = _T_1388 | io_exception; // @[CSR.scala 1021:17:freechips.rocketchip.system.DefaultRV32Config.fir@176695.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mprv = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_fs = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mstatus_mpp = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mstatus_spp = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_dcsr_prv = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_singleStepped = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_dcsr_ebreaku = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_debug = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_dcsr_cause = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  reg_dpc = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  reg_dscratch = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  reg_bp_0_control_dmode = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  reg_bp_0_control_action = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  reg_bp_0_control_tmatch = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  reg_bp_0_control_m = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  reg_bp_0_control_u = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  reg_bp_0_control_x = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  reg_bp_0_control_w = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  reg_bp_0_control_r = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  reg_bp_0_address = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  reg_pmp_0_cfg_l = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  reg_pmp_0_cfg_a = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  reg_pmp_0_cfg_x = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  reg_pmp_0_cfg_w = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  reg_pmp_0_cfg_r = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  reg_pmp_0_addr = _RAND_30[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  reg_pmp_1_cfg_l = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  reg_pmp_1_cfg_a = _RAND_32[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  reg_pmp_1_cfg_x = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  reg_pmp_1_cfg_w = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  reg_pmp_1_cfg_r = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  reg_pmp_1_addr = _RAND_36[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  reg_pmp_2_cfg_l = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  reg_pmp_2_cfg_a = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  reg_pmp_2_cfg_x = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  reg_pmp_2_cfg_w = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  reg_pmp_2_cfg_r = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  reg_pmp_2_addr = _RAND_42[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  reg_pmp_3_cfg_l = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  reg_pmp_3_cfg_a = _RAND_44[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  reg_pmp_3_cfg_x = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  reg_pmp_3_cfg_w = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  reg_pmp_3_cfg_r = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_pmp_3_addr = _RAND_48[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  reg_pmp_4_cfg_l = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  reg_pmp_4_cfg_a = _RAND_50[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  reg_pmp_4_cfg_x = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  reg_pmp_4_cfg_w = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  reg_pmp_4_cfg_r = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  reg_pmp_4_addr = _RAND_54[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  reg_pmp_5_cfg_l = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  reg_pmp_5_cfg_a = _RAND_56[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  reg_pmp_5_cfg_x = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  reg_pmp_5_cfg_w = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  reg_pmp_5_cfg_r = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  reg_pmp_5_addr = _RAND_60[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  reg_pmp_6_cfg_l = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  reg_pmp_6_cfg_a = _RAND_62[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  reg_pmp_6_cfg_x = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  reg_pmp_6_cfg_w = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  reg_pmp_6_cfg_r = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  reg_pmp_6_addr = _RAND_66[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  reg_pmp_7_cfg_l = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  reg_pmp_7_cfg_a = _RAND_68[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  reg_pmp_7_cfg_x = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  reg_pmp_7_cfg_w = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  reg_pmp_7_cfg_r = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  reg_pmp_7_addr = _RAND_72[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  reg_mie = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  reg_mepc = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  reg_mcause = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  reg_mtval = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  reg_mscratch = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  reg_mtvec = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  reg_mcounteren = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  reg_wfi = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  reg_fflags = _RAND_81[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  reg_frm = _RAND_82[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_87 = _RAND_83[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {2{`RANDOM}};
  _T_89 = _RAND_84[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_95 = _RAND_85[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  _T_97 = _RAND_86[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  reg_misa = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1387 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1743 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else begin
      if (_T_33) begin
        reg_mstatus_prv <= 2'h3;
      end else begin
        reg_mstatus_prv <= 2'h0;
      end
    end
    if (reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_604) begin
          reg_mstatus_mprv <= _T_4534;
        end
      end
    end
    if (reset) begin
      reg_mstatus_fs <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_604) begin
          if (_T_4555) begin
            reg_mstatus_fs <= 2'h3;
          end else begin
            reg_mstatus_fs <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_mpp <= 2'h3;
    end else begin
      if (csr_wen) begin
        if (_T_604) begin
          if (_T_4552) begin
            reg_mstatus_mpp <= 2'h3;
          end else begin
            reg_mstatus_mpp <= 2'h0;
          end
        end else begin
          if (insn_ret) begin
            if (_T_1729) begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  if (_T_1427) begin
                    reg_mstatus_mpp <= 2'h3;
                  end else begin
                    reg_mstatus_mpp <= 2'h0;
                  end
                end
              end
            end else begin
              reg_mstatus_mpp <= 2'h0;
            end
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (_T_1427) begin
                  reg_mstatus_mpp <= 2'h3;
                end else begin
                  reg_mstatus_mpp <= 2'h0;
                end
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_1729) begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (_T_1427) begin
                  reg_mstatus_mpp <= 2'h3;
                end else begin
                  reg_mstatus_mpp <= 2'h0;
                end
              end
            end
          end else begin
            reg_mstatus_mpp <= 2'h0;
          end
        end else begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (_T_1427) begin
                reg_mstatus_mpp <= 2'h3;
              end else begin
                reg_mstatus_mpp <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_spp <= 1'h0;
    end else begin
      reg_mstatus_spp <= _GEN_85[0];
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_604) begin
          reg_mstatus_mpie <= _T_4528;
        end else begin
          if (insn_ret) begin
            if (_T_1729) begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  reg_mstatus_mpie <= reg_mstatus_mie;
                end
              end
            end else begin
              reg_mstatus_mpie <= 1'h1;
            end
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_1729) begin
            if (exception) begin
              if (!(trapToDebug)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end else begin
            reg_mstatus_mpie <= 1'h1;
          end
        end else begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mpie <= reg_mstatus_mie;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_604) begin
          reg_mstatus_mie <= _T_4524;
        end else begin
          if (insn_ret) begin
            if (_T_1729) begin
              if (exception) begin
                reg_mstatus_mie <= _GEN_74;
              end
            end else begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end
          end else begin
            if (exception) begin
              reg_mstatus_mie <= _GEN_74;
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_1729) begin
            if (exception) begin
              reg_mstatus_mie <= _GEN_74;
            end
          end else begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end
        end else begin
          if (exception) begin
            reg_mstatus_mie <= _GEN_74;
          end
        end
      end
    end
    if (reset) begin
      reg_dcsr_prv <= 2'h3;
    end else begin
      if (csr_wen) begin
        if (_T_613) begin
          if (_T_4651) begin
            reg_dcsr_prv <= 2'h3;
          end else begin
            reg_dcsr_prv <= 2'h0;
          end
        end else begin
          if (exception) begin
            if (trapToDebug) begin
              if (_T_1423) begin
                reg_dcsr_prv <= _T_1429;
              end
            end
          end
        end
      end else begin
        if (exception) begin
          if (trapToDebug) begin
            if (_T_1423) begin
              reg_dcsr_prv <= _T_1429;
            end
          end
        end
      end
    end
    if (_T_277) begin
      reg_singleStepped <= 1'h0;
    end else begin
      reg_singleStepped <= _GEN_36;
    end
    if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_613) begin
          reg_dcsr_ebreakm <= _T_4647;
        end
      end
    end
    if (reset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_613) begin
          reg_dcsr_ebreaku <= _T_4644;
        end
      end
    end
    if (reset) begin
      reg_debug <= 1'h0;
    end else begin
      if (insn_ret) begin
        if (_T_1729) begin
          reg_debug <= 1'h0;
        end else begin
          if (exception) begin
            if (trapToDebug) begin
              reg_debug <= _GEN_38;
            end
          end
        end
      end else begin
        if (exception) begin
          if (trapToDebug) begin
            reg_debug <= _GEN_38;
          end
        end
      end
    end
    if (reset) begin
      reg_dcsr_cause <= 3'h0;
    end else begin
      if (exception) begin
        if (trapToDebug) begin
          if (_T_1423) begin
            if (reg_singleStepped) begin
              reg_dcsr_cause <= 3'h4;
            end else begin
              reg_dcsr_cause <= {{1'd0}, _T_1425};
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_613) begin
          reg_dcsr_step <= _T_4562;
        end
      end
    end
    if (csr_wen) begin
      if (_T_614) begin
        reg_dpc <= _T_4617;
      end else begin
        if (exception) begin
          if (trapToDebug) begin
            if (_T_1423) begin
              reg_dpc <= epc;
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (trapToDebug) begin
          if (_T_1423) begin
            reg_dpc <= epc;
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_615) begin
        reg_dscratch <= wdata;
      end
    end
    if (reset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4659) begin
          if (_T_601) begin
            reg_bp_0_control_dmode <= _T_4717;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_action <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4659) begin
          if (_T_601) begin
            reg_bp_0_control_action <= _GEN_158;
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_4659) begin
        if (_T_601) begin
          reg_bp_0_control_tmatch <= _T_4670;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4659) begin
        if (_T_601) begin
          reg_bp_0_control_m <= _T_4669;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4659) begin
        if (_T_601) begin
          reg_bp_0_control_u <= _T_4666;
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_x <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4659) begin
          if (_T_601) begin
            reg_bp_0_control_x <= _T_4562;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_w <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4659) begin
          if (_T_601) begin
            reg_bp_0_control_w <= _T_4664;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_r <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4659) begin
          if (_T_601) begin
            reg_bp_0_control_r <= _T_4663;
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_4659) begin
        if (_T_602) begin
          reg_bp_0_address <= wdata;
        end
      end
    end
    if (reset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4802) begin
          reg_pmp_0_cfg_l <= _T_4811;
        end
      end
    end
    if (reset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4802) begin
          reg_pmp_0_cfg_a <= _T_4809;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4802) begin
        reg_pmp_0_cfg_x <= _T_4808;
      end
    end
    if (csr_wen) begin
      if (_T_4802) begin
        reg_pmp_0_cfg_w <= _T_4812;
      end
    end
    if (csr_wen) begin
      if (_T_4802) begin
        reg_pmp_0_cfg_r <= _T_4806;
      end
    end
    reg_pmp_0_addr <= _GEN_353[29:0];
    if (reset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4822) begin
          reg_pmp_1_cfg_l <= _T_4831;
        end
      end
    end
    if (reset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4822) begin
          reg_pmp_1_cfg_a <= _T_4829;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4822) begin
        reg_pmp_1_cfg_x <= _T_4828;
      end
    end
    if (csr_wen) begin
      if (_T_4822) begin
        reg_pmp_1_cfg_w <= _T_4832;
      end
    end
    if (csr_wen) begin
      if (_T_4822) begin
        reg_pmp_1_cfg_r <= _T_4826;
      end
    end
    reg_pmp_1_addr <= _GEN_360[29:0];
    if (reset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4842) begin
          reg_pmp_2_cfg_l <= _T_4851;
        end
      end
    end
    if (reset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4842) begin
          reg_pmp_2_cfg_a <= _T_4849;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4842) begin
        reg_pmp_2_cfg_x <= _T_4848;
      end
    end
    if (csr_wen) begin
      if (_T_4842) begin
        reg_pmp_2_cfg_w <= _T_4852;
      end
    end
    if (csr_wen) begin
      if (_T_4842) begin
        reg_pmp_2_cfg_r <= _T_4846;
      end
    end
    reg_pmp_2_addr <= _GEN_367[29:0];
    if (reset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4862) begin
          reg_pmp_3_cfg_l <= _T_4871;
        end
      end
    end
    if (reset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4862) begin
          reg_pmp_3_cfg_a <= _T_4869;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4862) begin
        reg_pmp_3_cfg_x <= _T_4868;
      end
    end
    if (csr_wen) begin
      if (_T_4862) begin
        reg_pmp_3_cfg_w <= _T_4872;
      end
    end
    if (csr_wen) begin
      if (_T_4862) begin
        reg_pmp_3_cfg_r <= _T_4866;
      end
    end
    reg_pmp_3_addr <= _GEN_374[29:0];
    if (reset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4882) begin
          reg_pmp_4_cfg_l <= _T_4811;
        end
      end
    end
    if (reset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4882) begin
          reg_pmp_4_cfg_a <= _T_4809;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4882) begin
        reg_pmp_4_cfg_x <= _T_4808;
      end
    end
    if (csr_wen) begin
      if (_T_4882) begin
        reg_pmp_4_cfg_w <= _T_4812;
      end
    end
    if (csr_wen) begin
      if (_T_4882) begin
        reg_pmp_4_cfg_r <= _T_4806;
      end
    end
    reg_pmp_4_addr <= _GEN_381[29:0];
    if (reset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4902) begin
          reg_pmp_5_cfg_l <= _T_4831;
        end
      end
    end
    if (reset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4902) begin
          reg_pmp_5_cfg_a <= _T_4829;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4902) begin
        reg_pmp_5_cfg_x <= _T_4828;
      end
    end
    if (csr_wen) begin
      if (_T_4902) begin
        reg_pmp_5_cfg_w <= _T_4832;
      end
    end
    if (csr_wen) begin
      if (_T_4902) begin
        reg_pmp_5_cfg_r <= _T_4826;
      end
    end
    reg_pmp_5_addr <= _GEN_388[29:0];
    if (reset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4922) begin
          reg_pmp_6_cfg_l <= _T_4851;
        end
      end
    end
    if (reset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4922) begin
          reg_pmp_6_cfg_a <= _T_4849;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4922) begin
        reg_pmp_6_cfg_x <= _T_4848;
      end
    end
    if (csr_wen) begin
      if (_T_4922) begin
        reg_pmp_6_cfg_w <= _T_4852;
      end
    end
    if (csr_wen) begin
      if (_T_4922) begin
        reg_pmp_6_cfg_r <= _T_4846;
      end
    end
    reg_pmp_6_addr <= _GEN_395[29:0];
    if (reset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4942) begin
          reg_pmp_7_cfg_l <= _T_4871;
        end
      end
    end
    if (reset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_4942) begin
          reg_pmp_7_cfg_a <= _T_4869;
        end
      end
    end
    if (csr_wen) begin
      if (_T_4942) begin
        reg_pmp_7_cfg_x <= _T_4868;
      end
    end
    if (csr_wen) begin
      if (_T_4942) begin
        reg_pmp_7_cfg_w <= _T_4872;
      end
    end
    if (csr_wen) begin
      if (_T_4942) begin
        reg_pmp_7_cfg_r <= _T_4866;
      end
    end
    reg_pmp_7_addr <= _GEN_402[29:0];
    if (csr_wen) begin
      if (_T_607) begin
        reg_mie <= _T_4614;
      end
    end
    if (csr_wen) begin
      if (_T_609) begin
        reg_mepc <= _T_4617;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            reg_mepc <= epc;
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          reg_mepc <= epc;
        end
      end
    end
    if (csr_wen) begin
      if (_T_611) begin
        reg_mcause <= _T_4618;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (insn_call) begin
              reg_mcause <= {{28'd0}, _T_1334};
            end else begin
              if (insn_break) begin
                reg_mcause <= 32'h3;
              end else begin
                reg_mcause <= io_cause;
              end
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          if (insn_call) begin
            reg_mcause <= {{28'd0}, _T_1334};
          end else begin
            if (insn_break) begin
              reg_mcause <= 32'h3;
            end else begin
              reg_mcause <= io_cause;
            end
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_610) begin
        reg_mtval <= wdata;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            reg_mtval <= io_tval;
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          reg_mtval <= io_tval;
        end
      end
    end
    if (csr_wen) begin
      if (_T_608) begin
        reg_mscratch <= wdata;
      end
    end
    if (reset) begin
      reg_mtvec <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_605) begin
          reg_mtvec <= wdata;
        end
      end
    end
    if (csr_wen) begin
      if (_T_766) begin
        reg_mcounteren <= wdata;
      end
    end
    reg_fflags <= _GEN_305[4:0];
    reg_frm <= _GEN_306[2:0];
    if (reset) begin
      _T_87 <= 6'h0;
    end else begin
      _T_87 <= _GEN_302[5:0];
    end
    if (reset) begin
      _T_89 <= 58'h0;
    end else begin
      if (csr_wen) begin
        if (_T_770) begin
          _T_89 <= _T_4633;
        end else begin
          if (_T_620) begin
            _T_89 <= _T_4629;
          end else begin
            if (_T_90) begin
              _T_89 <= _T_92;
            end
          end
        end
      end else begin
        if (_T_90) begin
          _T_89 <= _T_92;
        end
      end
    end
    if (reset) begin
      reg_misa <= 32'h40901125;
    end else begin
      if (csr_wen) begin
        if (_T_603) begin
          if (_T_4563) begin
            reg_misa <= _T_4572;
          end
        end
      end
    end
    if (_T_1385) begin
      _T_1387 <= reg_mstatus_mpp;
    end else begin
      _T_1387 <= reg_mstatus_prv;
    end
    if (reset) begin
      _T_1743 <= 1'h0;
    end else begin
      _T_1743 <= _GEN_117;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1398) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:659 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@171693.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1398) begin
          $fatal; // @[CSR.scala 659:9:freechips.rocketchip.system.DefaultRV32Config.fir@171694.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1420) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:667 assert(!reg_singleStepped || io.retire === UInt(0))\n"); // @[CSR.scala 667:9:freechips.rocketchip.system.DefaultRV32Config.fir@171735.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1420) begin
          $fatal; // @[CSR.scala 667:9:freechips.rocketchip.system.DefaultRV32Config.fir@171736.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge io_ungated_clock) begin
    if (reset) begin
      reg_wfi <= 1'h0;
    end else begin
      if (_T_1405) begin
        reg_wfi <= 1'h0;
      end else begin
        reg_wfi <= _GEN_34;
      end
    end
    if (reset) begin
      _T_95 <= 6'h0;
    end else begin
      _T_95 <= _GEN_300[5:0];
    end
    if (reset) begin
      _T_97 <= 58'h0;
    end else begin
      if (csr_wen) begin
        if (_T_769) begin
          _T_97 <= _T_4626;
        end else begin
          if (_T_619) begin
            _T_97 <= _T_4622;
          end else begin
            if (_T_98) begin
              _T_97 <= _T_100;
            end
          end
        end
      end else begin
        if (_T_98) begin
          _T_97 <= _T_100;
        end
      end
    end
  end
endmodule
`endif // __CSRFile
