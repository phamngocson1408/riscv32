
module TLROM( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195903.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195904.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195905.4]
  output        auto_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input         auto_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input  [2:0]  auto_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input  [2:0]  auto_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input  [1:0]  auto_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input  [9:0]  auto_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input  [16:0] auto_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input  [3:0]  auto_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input         auto_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  input         auto_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  output        auto_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  output [1:0]  auto_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  output [9:0]  auto_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
  output [31:0] auto_in_d_bits_data // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195906.4]
);
  wire  TLMonitor_clock; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [1:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [9:0] TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [16:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [3:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire  TLMonitor_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [1:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [9:0] TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
  wire [9:0] index; // @[BootROM.scala 50:34:freechips.rocketchip.system.DefaultRV32Config.fir@196965.4]
  wire [3:0] high; // @[BootROM.scala 51:68:freechips.rocketchip.system.DefaultRV32Config.fir@196966.4]
  wire  _T; // @[BootROM.scala 52:53:freechips.rocketchip.system.DefaultRV32Config.fir@196967.4]
  wire [31:0] _GEN_1; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_2; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_3; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_4; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_5; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_6; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_7; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_8; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_9; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_10; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_11; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_12; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_13; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_14; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_15; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_16; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_17; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_18; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_19; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_20; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_21; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_22; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_23; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_24; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_25; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_26; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_27; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_28; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_29; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_30; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_31; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_32; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_33; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_34; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_35; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_36; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_37; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_38; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_39; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_40; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_41; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_42; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_43; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_44; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_45; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_46; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_47; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_48; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_49; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_50; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_51; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_52; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_53; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_54; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_55; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_56; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_57; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_58; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_59; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_60; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_61; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_62; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_63; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_64; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_65; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_66; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_67; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_68; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_69; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_70; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_71; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_72; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_73; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_74; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_75; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_76; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_77; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_78; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_79; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_80; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_81; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_82; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_83; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_84; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_85; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_86; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_87; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_88; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_89; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_90; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_91; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_92; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_93; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_94; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_95; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_96; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_97; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_98; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_99; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_100; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_101; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_102; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_103; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_104; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_105; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_106; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_107; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_108; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_109; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_110; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_111; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_112; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_113; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_114; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_115; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_116; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_117; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_118; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_119; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_120; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_121; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_122; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_123; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_124; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_125; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_126; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_127; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_128; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_129; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_130; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_131; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_132; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_133; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_134; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_135; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_136; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_137; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_138; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_139; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_140; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_141; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_142; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_143; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_144; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_145; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_146; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_147; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_148; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_149; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_150; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_151; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_152; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_153; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_154; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_155; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_156; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_157; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_158; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_159; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_160; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_161; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_162; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_163; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_164; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_165; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_166; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_167; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_168; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_169; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_170; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_171; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_172; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_173; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_174; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_175; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_176; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_177; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_178; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_179; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_180; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_181; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_182; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_183; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_184; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_185; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_186; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_187; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_188; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_189; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_190; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_191; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_192; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_193; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_194; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_195; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_196; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_197; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_198; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_199; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_200; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_201; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_202; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_203; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_204; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_205; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_206; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_207; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_208; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_209; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_210; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_211; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_212; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_213; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_214; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_215; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_216; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_217; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_218; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_219; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_220; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_221; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_222; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_223; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_224; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_225; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_226; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_227; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_228; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_229; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_230; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_231; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_232; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_233; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_234; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_235; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_236; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_237; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_238; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_239; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_240; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_241; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_242; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_243; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_244; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_245; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_246; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_247; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_248; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_249; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_250; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_251; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_252; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_253; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_254; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_255; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_256; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_257; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_258; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_259; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_260; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_261; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_262; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_263; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_264; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_265; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_266; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_267; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_268; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_269; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_270; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_271; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_272; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_273; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_274; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_275; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_276; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_277; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_278; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_279; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_280; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_281; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_282; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_283; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_284; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_285; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_286; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_287; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_288; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_289; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_290; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_291; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_292; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_293; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_294; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_295; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_296; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_297; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_298; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_299; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_300; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_301; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_302; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_303; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_304; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_305; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_306; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_307; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_308; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_309; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_310; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_311; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_312; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_313; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_314; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_315; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_316; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_317; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_318; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_319; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_320; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_321; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_322; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_323; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_324; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_325; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_326; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_327; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_328; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_329; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_330; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_331; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_332; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_333; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_334; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_335; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_336; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_337; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_338; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_339; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_340; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_341; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_342; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_343; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_344; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_345; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_346; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_347; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_348; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_349; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_350; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_351; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_352; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_353; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_354; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_355; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_356; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_357; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_358; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_359; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_360; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_361; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_362; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_363; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_364; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_365; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_366; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_367; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_368; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_369; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_370; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_371; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_372; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_373; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_374; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_375; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_376; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_377; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_378; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_379; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_380; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_381; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_382; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_383; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_384; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_385; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_386; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_387; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_388; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_389; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_390; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_391; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_392; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_393; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_394; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_395; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_396; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_397; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_398; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_399; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_400; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_401; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_402; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_403; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_404; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_405; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_406; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_407; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_408; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_409; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_410; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_411; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_412; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_413; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_414; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_415; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_416; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_417; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_418; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_419; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_420; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_421; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_422; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_423; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_424; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_425; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_426; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_427; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_428; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_429; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_430; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_431; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_432; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_433; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_434; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_435; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_436; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_437; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_438; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_439; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_440; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_441; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_442; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_443; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_444; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_445; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_446; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_447; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_448; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_449; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_450; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_451; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_452; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_453; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_454; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_455; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_456; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_457; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_458; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_459; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_460; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_461; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_462; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_463; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_464; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_465; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_466; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_467; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_468; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_469; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_470; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_471; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_472; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_473; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_474; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_475; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_476; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_477; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_478; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_479; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_480; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_481; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_482; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_483; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_484; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_485; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_486; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_487; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_488; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_489; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_490; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_491; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_492; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_493; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_494; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_495; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_496; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_497; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_498; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_499; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_500; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_501; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_502; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_503; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_504; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_505; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_506; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_507; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_508; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_509; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_510; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_511; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_512; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_513; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_514; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_515; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_516; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_517; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_518; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_519; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_520; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_521; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_522; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_523; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_524; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_525; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_526; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_527; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_528; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_529; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_530; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_531; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_532; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_533; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_534; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_535; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_536; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_537; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_538; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_539; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_540; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_541; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_542; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_543; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_544; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_545; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_546; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_547; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_548; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_549; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_550; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_551; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_552; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_553; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_554; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_555; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_556; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_557; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_558; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_559; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_560; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_561; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_562; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_563; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_564; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_565; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_566; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_567; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_568; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_569; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_570; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_571; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_572; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_573; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_574; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_575; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_576; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_577; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_578; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_579; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_580; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_581; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_582; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_583; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_584; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_585; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_586; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_587; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_588; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_589; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_590; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_591; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_592; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_593; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_594; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_595; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_596; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_597; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_598; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_599; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_600; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_601; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_602; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_603; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_604; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_605; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_606; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_607; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_608; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_609; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_610; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_611; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_612; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_613; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_614; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_615; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_616; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_617; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_618; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_619; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_620; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_621; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_622; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_623; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_624; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_625; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_626; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_627; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_628; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_629; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_630; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_631; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_632; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_633; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_634; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_635; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_636; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_637; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_638; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_639; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_640; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_641; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_642; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_643; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_644; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_645; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_646; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_647; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_648; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_649; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_650; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_651; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_652; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_653; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_654; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_655; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_656; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_657; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_658; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_659; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_660; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_661; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_662; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_663; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_664; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_665; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_666; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_667; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_668; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_669; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_670; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_671; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_672; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_673; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_674; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_675; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_676; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_677; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_678; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_679; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_680; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_681; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_682; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_683; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_684; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_685; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_686; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_687; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_688; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_689; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_690; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_691; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_692; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_693; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_694; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_695; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_696; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_697; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_698; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_699; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_700; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_701; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_702; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_703; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_704; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_705; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_706; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_707; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_708; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_709; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_710; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_711; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_712; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_713; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_714; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_715; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_716; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_717; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_718; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_719; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_720; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_721; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_722; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_723; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_724; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_725; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_726; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_727; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_728; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_729; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_730; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_731; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_732; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_733; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_734; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_735; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_736; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_737; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_738; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_739; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_740; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_741; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_742; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_743; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_744; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_745; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_746; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_747; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_748; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_749; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_750; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_751; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_752; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_753; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_754; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_755; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_756; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_757; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_758; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_759; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_760; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_761; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_762; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_763; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_764; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_765; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_766; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_767; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_768; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_769; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_770; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_771; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_772; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_773; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_774; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_775; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_776; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_777; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_778; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_779; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_780; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_781; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_782; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_783; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_784; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_785; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_786; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_787; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_788; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_789; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_790; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_791; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_792; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_793; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_794; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_795; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_796; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_797; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_798; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_799; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_800; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_801; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_802; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_803; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_804; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_805; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_806; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_807; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_808; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_809; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_810; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_811; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_812; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_813; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_814; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_815; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_816; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_817; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_818; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_819; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_820; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_821; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_822; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_823; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_824; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_825; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_826; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_827; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_828; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_829; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_830; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_831; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_832; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_833; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_834; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_835; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_836; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_837; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_838; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_839; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_840; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_841; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_842; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_843; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_844; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_845; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_846; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_847; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_848; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_849; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_850; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_851; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_852; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_853; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_854; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_855; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_856; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_857; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_858; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_859; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_860; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_861; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_862; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_863; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_864; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_865; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_866; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_867; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_868; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_869; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_870; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_871; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_872; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_873; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_874; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_875; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_876; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_877; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_878; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_879; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_880; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_881; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_882; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_883; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_884; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_885; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_886; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_887; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_888; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_889; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_890; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_891; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_892; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_893; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_894; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_895; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_896; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_897; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_898; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_899; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_900; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_901; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_902; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_903; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_904; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_905; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_906; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_907; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_908; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_909; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_910; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_911; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_912; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_913; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_914; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_915; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_916; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_917; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_918; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_919; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_920; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_921; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_922; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_923; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_924; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_925; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_926; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_927; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_928; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_929; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_930; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_931; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_932; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_933; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_934; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_935; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_936; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_937; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_938; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_939; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_940; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_941; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_942; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_943; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_944; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_945; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_946; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_947; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_948; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_949; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_950; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_951; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_952; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_953; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_954; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_955; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_956; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_957; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_958; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_959; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_960; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_961; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_962; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_963; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_964; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_965; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_966; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_967; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_968; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_969; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_970; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_971; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_972; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_973; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_974; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_975; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_976; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_977; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_978; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_979; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_980; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_981; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_982; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_983; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_984; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_985; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_986; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_987; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_988; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_989; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_990; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_991; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_992; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_993; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_994; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_995; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_996; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_997; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_998; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_999; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1000; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1001; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1002; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1003; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1004; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1005; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1006; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1007; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1008; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1009; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1010; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1011; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1012; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1013; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1014; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1015; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1016; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1017; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1018; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1019; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1020; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1021; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1022; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  wire [31:0] _GEN_1023; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  TLMonitor_45 TLMonitor ( // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultRV32Config.fir@195913.4]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source)
  );
  assign index = auto_in_a_bits_address[11:2]; // @[BootROM.scala 50:34:freechips.rocketchip.system.DefaultRV32Config.fir@196965.4]
  assign high = auto_in_a_bits_address[15:12]; // @[BootROM.scala 51:68:freechips.rocketchip.system.DefaultRV32Config.fir@196966.4]
  assign _T = high != 4'h0; // @[BootROM.scala 52:53:freechips.rocketchip.system.DefaultRV32Config.fir@196967.4]
  assign _GEN_1 = 10'h1 == index ? 32'h1f41413 : 32'h10041b; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_2 = 10'h2 == index ? 32'hf1402573 : _GEN_1; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_3 = 10'h3 == index ? 32'h597 : _GEN_2; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_4 = 10'h4 == index ? 32'h7458593 : _GEN_3; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_5 = 10'h5 == index ? 32'h8402 : _GEN_4; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_6 = 10'h6 == index ? 32'h0 : _GEN_5; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_7 = 10'h7 == index ? 32'h0 : _GEN_6; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_8 = 10'h8 == index ? 32'h0 : _GEN_7; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_9 = 10'h9 == index ? 32'h0 : _GEN_8; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_10 = 10'ha == index ? 32'h0 : _GEN_9; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_11 = 10'hb == index ? 32'h0 : _GEN_10; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_12 = 10'hc == index ? 32'h0 : _GEN_11; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_13 = 10'hd == index ? 32'h0 : _GEN_12; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_14 = 10'he == index ? 32'h0 : _GEN_13; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_15 = 10'hf == index ? 32'h0 : _GEN_14; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_16 = 10'h10 == index ? 32'hf1402573 : _GEN_15; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_17 = 10'h11 == index ? 32'h597 : _GEN_16; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_18 = 10'h12 == index ? 32'h3c58593 : _GEN_17; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_19 = 10'h13 == index ? 32'h8137 : _GEN_18; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_20 = 10'h14 == index ? 32'h11011b : _GEN_19; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_21 = 10'h15 == index ? 32'h1011113 : _GEN_20; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_22 = 10'h16 == index ? 32'h10061b : _GEN_21; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_23 = 10'h17 == index ? 32'h1f61613 : _GEN_22; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_24 = 10'h18 == index ? 32'ha0018602 : _GEN_23; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_25 = 10'h19 == index ? 32'h0 : _GEN_24; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_26 = 10'h1a == index ? 32'h0 : _GEN_25; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_27 = 10'h1b == index ? 32'h0 : _GEN_26; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_28 = 10'h1c == index ? 32'h0 : _GEN_27; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_29 = 10'h1d == index ? 32'h0 : _GEN_28; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_30 = 10'h1e == index ? 32'h0 : _GEN_29; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_31 = 10'h1f == index ? 32'h0 : _GEN_30; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_32 = 10'h20 == index ? 32'hedfe0dd0 : _GEN_31; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_33 = 10'h21 == index ? 32'hc0080000 : _GEN_32; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_34 = 10'h22 == index ? 32'h38000000 : _GEN_33; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_35 = 10'h23 == index ? 32'hdc060000 : _GEN_34; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_36 = 10'h24 == index ? 32'h28000000 : _GEN_35; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_37 = 10'h25 == index ? 32'h11000000 : _GEN_36; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_38 = 10'h26 == index ? 32'h10000000 : _GEN_37; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_39 = 10'h27 == index ? 32'h0 : _GEN_38; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_40 = 10'h28 == index ? 32'he4010000 : _GEN_39; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_41 = 10'h29 == index ? 32'ha4060000 : _GEN_40; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_42 = 10'h2a == index ? 32'h0 : _GEN_41; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_43 = 10'h2b == index ? 32'h0 : _GEN_42; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_44 = 10'h2c == index ? 32'h0 : _GEN_43; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_45 = 10'h2d == index ? 32'h0 : _GEN_44; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_46 = 10'h2e == index ? 32'h1000000 : _GEN_45; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_47 = 10'h2f == index ? 32'h0 : _GEN_46; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_48 = 10'h30 == index ? 32'h3000000 : _GEN_47; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_49 = 10'h31 == index ? 32'h4000000 : _GEN_48; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_50 = 10'h32 == index ? 32'h0 : _GEN_49; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_51 = 10'h33 == index ? 32'h1000000 : _GEN_50; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_52 = 10'h34 == index ? 32'h3000000 : _GEN_51; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_53 = 10'h35 == index ? 32'h4000000 : _GEN_52; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_54 = 10'h36 == index ? 32'hf000000 : _GEN_53; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_55 = 10'h37 == index ? 32'h1000000 : _GEN_54; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_56 = 10'h38 == index ? 32'h3000000 : _GEN_55; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_57 = 10'h39 == index ? 32'h21000000 : _GEN_56; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_58 = 10'h3a == index ? 32'h1b000000 : _GEN_57; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_59 = 10'h3b == index ? 32'h65657266 : _GEN_58; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_60 = 10'h3c == index ? 32'h70696863 : _GEN_59; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_61 = 10'h3d == index ? 32'h6f722c73 : _GEN_60; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_62 = 10'h3e == index ? 32'h74656b63 : _GEN_61; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_63 = 10'h3f == index ? 32'h70696863 : _GEN_62; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_64 = 10'h40 == index ? 32'h6b6e752d : _GEN_63; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_65 = 10'h41 == index ? 32'h6e776f6e : _GEN_64; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_66 = 10'h42 == index ? 32'h7665642d : _GEN_65; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_67 = 10'h43 == index ? 32'h0 : _GEN_66; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_68 = 10'h44 == index ? 32'h3000000 : _GEN_67; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_69 = 10'h45 == index ? 32'h1d000000 : _GEN_68; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_70 = 10'h46 == index ? 32'h26000000 : _GEN_69; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_71 = 10'h47 == index ? 32'h65657266 : _GEN_70; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_72 = 10'h48 == index ? 32'h70696863 : _GEN_71; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_73 = 10'h49 == index ? 32'h6f722c73 : _GEN_72; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_74 = 10'h4a == index ? 32'h74656b63 : _GEN_73; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_75 = 10'h4b == index ? 32'h70696863 : _GEN_74; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_76 = 10'h4c == index ? 32'h6b6e752d : _GEN_75; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_77 = 10'h4d == index ? 32'h6e776f6e : _GEN_76; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_78 = 10'h4e == index ? 32'h0 : _GEN_77; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_79 = 10'h4f == index ? 32'h1000000 : _GEN_78; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_80 = 10'h50 == index ? 32'h73757063 : _GEN_79; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_81 = 10'h51 == index ? 32'h0 : _GEN_80; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_82 = 10'h52 == index ? 32'h3000000 : _GEN_81; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_83 = 10'h53 == index ? 32'h4000000 : _GEN_82; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_84 = 10'h54 == index ? 32'h0 : _GEN_83; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_85 = 10'h55 == index ? 32'h1000000 : _GEN_84; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_86 = 10'h56 == index ? 32'h3000000 : _GEN_85; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_87 = 10'h57 == index ? 32'h4000000 : _GEN_86; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_88 = 10'h58 == index ? 32'hf000000 : _GEN_87; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_89 = 10'h59 == index ? 32'h0 : _GEN_88; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_90 = 10'h5a == index ? 32'h1000000 : _GEN_89; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_91 = 10'h5b == index ? 32'h40757063 : _GEN_90; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_92 = 10'h5c == index ? 32'h30 : _GEN_91; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_93 = 10'h5d == index ? 32'h3000000 : _GEN_92; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_94 = 10'h5e == index ? 32'h4000000 : _GEN_93; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_95 = 10'h5f == index ? 32'h2c000000 : _GEN_94; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_96 = 10'h60 == index ? 32'h0 : _GEN_95; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_97 = 10'h61 == index ? 32'h3000000 : _GEN_96; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_98 = 10'h62 == index ? 32'h15000000 : _GEN_97; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_99 = 10'h63 == index ? 32'h1b000000 : _GEN_98; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_100 = 10'h64 == index ? 32'h69666973 : _GEN_99; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_101 = 10'h65 == index ? 32'h722c6576 : _GEN_100; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_102 = 10'h66 == index ? 32'h656b636f : _GEN_101; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_103 = 10'h67 == index ? 32'h72003074 : _GEN_102; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_104 = 10'h68 == index ? 32'h76637369 : _GEN_103; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_105 = 10'h69 == index ? 32'h0 : _GEN_104; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_106 = 10'h6a == index ? 32'h3000000 : _GEN_105; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_107 = 10'h6b == index ? 32'h4000000 : _GEN_106; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_108 = 10'h6c == index ? 32'h3c000000 : _GEN_107; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_109 = 10'h6d == index ? 32'h40000000 : _GEN_108; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_110 = 10'h6e == index ? 32'h3000000 : _GEN_109; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_111 = 10'h6f == index ? 32'h4000000 : _GEN_110; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_112 = 10'h70 == index ? 32'h4f000000 : _GEN_111; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_113 = 10'h71 == index ? 32'h40000000 : _GEN_112; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_114 = 10'h72 == index ? 32'h3000000 : _GEN_113; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_115 = 10'h73 == index ? 32'h4000000 : _GEN_114; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_116 = 10'h74 == index ? 32'h5c000000 : _GEN_115; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_117 = 10'h75 == index ? 32'h400000 : _GEN_116; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_118 = 10'h76 == index ? 32'h3000000 : _GEN_117; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_119 = 10'h77 == index ? 32'h4000000 : _GEN_118; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_120 = 10'h78 == index ? 32'h69000000 : _GEN_119; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_121 = 10'h79 == index ? 32'h1000000 : _GEN_120; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_122 = 10'h7a == index ? 32'h3000000 : _GEN_121; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_123 = 10'h7b == index ? 32'h4000000 : _GEN_122; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_124 = 10'h7c == index ? 32'h74000000 : _GEN_123; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_125 = 10'h7d == index ? 32'h20000000 : _GEN_124; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_126 = 10'h7e == index ? 32'h3000000 : _GEN_125; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_127 = 10'h7f == index ? 32'h4000000 : _GEN_126; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_128 = 10'h80 == index ? 32'h7f000000 : _GEN_127; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_129 = 10'h81 == index ? 32'h757063 : _GEN_128; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_130 = 10'h82 == index ? 32'h3000000 : _GEN_129; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_131 = 10'h83 == index ? 32'h4000000 : _GEN_130; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_132 = 10'h84 == index ? 32'h8b000000 : _GEN_131; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_133 = 10'h85 == index ? 32'h1000000 : _GEN_132; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_134 = 10'h86 == index ? 32'h3000000 : _GEN_133; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_135 = 10'h87 == index ? 32'h4000000 : _GEN_134; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_136 = 10'h88 == index ? 32'haa000000 : _GEN_135; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_137 = 10'h89 == index ? 32'h40000000 : _GEN_136; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_138 = 10'h8a == index ? 32'h3000000 : _GEN_137; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_139 = 10'h8b == index ? 32'h4000000 : _GEN_138; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_140 = 10'h8c == index ? 32'hbd000000 : _GEN_139; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_141 = 10'h8d == index ? 32'h40000000 : _GEN_140; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_142 = 10'h8e == index ? 32'h3000000 : _GEN_141; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_143 = 10'h8f == index ? 32'h4000000 : _GEN_142; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_144 = 10'h90 == index ? 32'hca000000 : _GEN_143; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_145 = 10'h91 == index ? 32'h400000 : _GEN_144; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_146 = 10'h92 == index ? 32'h3000000 : _GEN_145; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_147 = 10'h93 == index ? 32'h4000000 : _GEN_146; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_148 = 10'h94 == index ? 32'hd7000000 : _GEN_147; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_149 = 10'h95 == index ? 32'h1000000 : _GEN_148; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_150 = 10'h96 == index ? 32'h3000000 : _GEN_149; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_151 = 10'h97 == index ? 32'h4000000 : _GEN_150; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_152 = 10'h98 == index ? 32'he2000000 : _GEN_151; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_153 = 10'h99 == index ? 32'h20000000 : _GEN_152; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_154 = 10'h9a == index ? 32'h3000000 : _GEN_153; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_155 = 10'h9b == index ? 32'hb000000 : _GEN_154; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_156 = 10'h9c == index ? 32'hed000000 : _GEN_155; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_157 = 10'h9d == index ? 32'h63736972 : _GEN_156; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_158 = 10'h9e == index ? 32'h76732c76 : _GEN_157; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_159 = 10'h9f == index ? 32'h3233 : _GEN_158; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_160 = 10'ha0 == index ? 32'h3000000 : _GEN_159; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_161 = 10'ha1 == index ? 32'h4000000 : _GEN_160; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_162 = 10'ha2 == index ? 32'hf6000000 : _GEN_161; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_163 = 10'ha3 == index ? 32'h1000000 : _GEN_162; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_164 = 10'ha4 == index ? 32'h3000000 : _GEN_163; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_165 = 10'ha5 == index ? 32'h4000000 : _GEN_164; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_166 = 10'ha6 == index ? 32'h7010000 : _GEN_165; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_167 = 10'ha7 == index ? 32'h0 : _GEN_166; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_168 = 10'ha8 == index ? 32'h3000000 : _GEN_167; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_169 = 10'ha9 == index ? 32'ha000000 : _GEN_168; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_170 = 10'haa == index ? 32'hb010000 : _GEN_169; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_171 = 10'hab == index ? 32'h32337672 : _GEN_170; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_172 = 10'hac == index ? 32'h66616d69 : _GEN_171; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_173 = 10'had == index ? 32'h63 : _GEN_172; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_174 = 10'hae == index ? 32'h3000000 : _GEN_173; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_175 = 10'haf == index ? 32'h4000000 : _GEN_174; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_176 = 10'hb0 == index ? 32'h15010000 : _GEN_175; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_177 = 10'hb1 == index ? 32'h8000000 : _GEN_176; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_178 = 10'hb2 == index ? 32'h3000000 : _GEN_177; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_179 = 10'hb3 == index ? 32'h5000000 : _GEN_178; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_180 = 10'hb4 == index ? 32'h26010000 : _GEN_179; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_181 = 10'hb5 == index ? 32'h79616b6f : _GEN_180; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_182 = 10'hb6 == index ? 32'h0 : _GEN_181; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_183 = 10'hb7 == index ? 32'h3000000 : _GEN_182; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_184 = 10'hb8 == index ? 32'h4000000 : _GEN_183; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_185 = 10'hb9 == index ? 32'h2d010000 : _GEN_184; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_186 = 10'hba == index ? 32'h40420f00 : _GEN_185; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_187 = 10'hbb == index ? 32'h3000000 : _GEN_186; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_188 = 10'hbc == index ? 32'h0 : _GEN_187; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_189 = 10'hbd == index ? 32'h40010000 : _GEN_188; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_190 = 10'hbe == index ? 32'h1000000 : _GEN_189; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_191 = 10'hbf == index ? 32'h65746e69 : _GEN_190; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_192 = 10'hc0 == index ? 32'h70757272 : _GEN_191; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_193 = 10'hc1 == index ? 32'h6f632d74 : _GEN_192; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_194 = 10'hc2 == index ? 32'h6f72746e : _GEN_193; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_195 = 10'hc3 == index ? 32'h72656c6c : _GEN_194; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_196 = 10'hc4 == index ? 32'h0 : _GEN_195; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_197 = 10'hc5 == index ? 32'h3000000 : _GEN_196; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_198 = 10'hc6 == index ? 32'h4000000 : _GEN_197; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_199 = 10'hc7 == index ? 32'h4a010000 : _GEN_198; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_200 = 10'hc8 == index ? 32'h1000000 : _GEN_199; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_201 = 10'hc9 == index ? 32'h3000000 : _GEN_200; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_202 = 10'hca == index ? 32'hf000000 : _GEN_201; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_203 = 10'hcb == index ? 32'h1b000000 : _GEN_202; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_204 = 10'hcc == index ? 32'h63736972 : _GEN_203; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_205 = 10'hcd == index ? 32'h70632c76 : _GEN_204; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_206 = 10'hce == index ? 32'h6e692d75 : _GEN_205; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_207 = 10'hcf == index ? 32'h6374 : _GEN_206; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_208 = 10'hd0 == index ? 32'h3000000 : _GEN_207; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_209 = 10'hd1 == index ? 32'h0 : _GEN_208; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_210 = 10'hd2 == index ? 32'h5b010000 : _GEN_209; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_211 = 10'hd3 == index ? 32'h3000000 : _GEN_210; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_212 = 10'hd4 == index ? 32'h4000000 : _GEN_211; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_213 = 10'hd5 == index ? 32'h70010000 : _GEN_212; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_214 = 10'hd6 == index ? 32'h2000000 : _GEN_213; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_215 = 10'hd7 == index ? 32'h2000000 : _GEN_214; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_216 = 10'hd8 == index ? 32'h2000000 : _GEN_215; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_217 = 10'hd9 == index ? 32'h2000000 : _GEN_216; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_218 = 10'hda == index ? 32'h1000000 : _GEN_217; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_219 = 10'hdb == index ? 32'h6f6d656d : _GEN_218; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_220 = 10'hdc == index ? 32'h38407972 : _GEN_219; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_221 = 10'hdd == index ? 32'h30303030 : _GEN_220; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_222 = 10'hde == index ? 32'h303030 : _GEN_221; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_223 = 10'hdf == index ? 32'h3000000 : _GEN_222; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_224 = 10'he0 == index ? 32'h7000000 : _GEN_223; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_225 = 10'he1 == index ? 32'h7f000000 : _GEN_224; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_226 = 10'he2 == index ? 32'h6f6d656d : _GEN_225; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_227 = 10'he3 == index ? 32'h7972 : _GEN_226; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_228 = 10'he4 == index ? 32'h3000000 : _GEN_227; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_229 = 10'he5 == index ? 32'h8000000 : _GEN_228; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_230 = 10'he6 == index ? 32'h7010000 : _GEN_229; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_231 = 10'he7 == index ? 32'h80 : _GEN_230; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_232 = 10'he8 == index ? 32'h10 : _GEN_231; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_233 = 10'he9 == index ? 32'h3000000 : _GEN_232; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_234 = 10'hea == index ? 32'h4000000 : _GEN_233; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_235 = 10'heb == index ? 32'h70010000 : _GEN_234; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_236 = 10'hec == index ? 32'h1000000 : _GEN_235; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_237 = 10'hed == index ? 32'h2000000 : _GEN_236; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_238 = 10'hee == index ? 32'h1000000 : _GEN_237; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_239 = 10'hef == index ? 32'h636f73 : _GEN_238; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_240 = 10'hf0 == index ? 32'h3000000 : _GEN_239; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_241 = 10'hf1 == index ? 32'h4000000 : _GEN_240; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_242 = 10'hf2 == index ? 32'h0 : _GEN_241; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_243 = 10'hf3 == index ? 32'h1000000 : _GEN_242; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_244 = 10'hf4 == index ? 32'h3000000 : _GEN_243; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_245 = 10'hf5 == index ? 32'h4000000 : _GEN_244; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_246 = 10'hf6 == index ? 32'hf000000 : _GEN_245; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_247 = 10'hf7 == index ? 32'h1000000 : _GEN_246; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_248 = 10'hf8 == index ? 32'h3000000 : _GEN_247; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_249 = 10'hf9 == index ? 32'h2c000000 : _GEN_248; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_250 = 10'hfa == index ? 32'h1b000000 : _GEN_249; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_251 = 10'hfb == index ? 32'h65657266 : _GEN_250; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_252 = 10'hfc == index ? 32'h70696863 : _GEN_251; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_253 = 10'hfd == index ? 32'h6f722c73 : _GEN_252; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_254 = 10'hfe == index ? 32'h74656b63 : _GEN_253; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_255 = 10'hff == index ? 32'h70696863 : _GEN_254; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_256 = 10'h100 == index ? 32'h6b6e752d : _GEN_255; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_257 = 10'h101 == index ? 32'h6e776f6e : _GEN_256; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_258 = 10'h102 == index ? 32'h636f732d : _GEN_257; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_259 = 10'h103 == index ? 32'h6d697300 : _GEN_258; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_260 = 10'h104 == index ? 32'h2d656c70 : _GEN_259; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_261 = 10'h105 == index ? 32'h737562 : _GEN_260; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_262 = 10'h106 == index ? 32'h3000000 : _GEN_261; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_263 = 10'h107 == index ? 32'h0 : _GEN_262; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_264 = 10'h108 == index ? 32'h78010000 : _GEN_263; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_265 = 10'h109 == index ? 32'h1000000 : _GEN_264; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_266 = 10'h10a == index ? 32'h6e696c63 : _GEN_265; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_267 = 10'h10b == index ? 32'h30324074 : _GEN_266; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_268 = 10'h10c == index ? 32'h30303030 : _GEN_267; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_269 = 10'h10d == index ? 32'h30 : _GEN_268; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_270 = 10'h10e == index ? 32'h3000000 : _GEN_269; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_271 = 10'h10f == index ? 32'hd000000 : _GEN_270; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_272 = 10'h110 == index ? 32'h1b000000 : _GEN_271; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_273 = 10'h111 == index ? 32'h63736972 : _GEN_272; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_274 = 10'h112 == index ? 32'h6c632c76 : _GEN_273; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_275 = 10'h113 == index ? 32'h30746e69 : _GEN_274; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_276 = 10'h114 == index ? 32'h0 : _GEN_275; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_277 = 10'h115 == index ? 32'h3000000 : _GEN_276; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_278 = 10'h116 == index ? 32'h10000000 : _GEN_277; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_279 = 10'h117 == index ? 32'h7f010000 : _GEN_278; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_280 = 10'h118 == index ? 32'h2000000 : _GEN_279; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_281 = 10'h119 == index ? 32'h3000000 : _GEN_280; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_282 = 10'h11a == index ? 32'h2000000 : _GEN_281; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_283 = 10'h11b == index ? 32'h7000000 : _GEN_282; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_284 = 10'h11c == index ? 32'h3000000 : _GEN_283; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_285 = 10'h11d == index ? 32'h8000000 : _GEN_284; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_286 = 10'h11e == index ? 32'h7010000 : _GEN_285; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_287 = 10'h11f == index ? 32'h2 : _GEN_286; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_288 = 10'h120 == index ? 32'h100 : _GEN_287; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_289 = 10'h121 == index ? 32'h3000000 : _GEN_288; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_290 = 10'h122 == index ? 32'h8000000 : _GEN_289; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_291 = 10'h123 == index ? 32'h93010000 : _GEN_290; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_292 = 10'h124 == index ? 32'h746e6f63 : _GEN_291; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_293 = 10'h125 == index ? 32'h6c6f72 : _GEN_292; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_294 = 10'h126 == index ? 32'h2000000 : _GEN_293; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_295 = 10'h127 == index ? 32'h1000000 : _GEN_294; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_296 = 10'h128 == index ? 32'h75626564 : _GEN_295; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_297 = 10'h129 == index ? 32'h6f632d67 : _GEN_296; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_298 = 10'h12a == index ? 32'h6f72746e : _GEN_297; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_299 = 10'h12b == index ? 32'h72656c6c : _GEN_298; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_300 = 10'h12c == index ? 32'h3040 : _GEN_299; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_301 = 10'h12d == index ? 32'h3000000 : _GEN_300; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_302 = 10'h12e == index ? 32'h21000000 : _GEN_301; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_303 = 10'h12f == index ? 32'h1b000000 : _GEN_302; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_304 = 10'h130 == index ? 32'h69666973 : _GEN_303; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_305 = 10'h131 == index ? 32'h642c6576 : _GEN_304; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_306 = 10'h132 == index ? 32'h67756265 : _GEN_305; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_307 = 10'h133 == index ? 32'h3331302d : _GEN_306; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_308 = 10'h134 == index ? 32'h73697200 : _GEN_307; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_309 = 10'h135 == index ? 32'h642c7663 : _GEN_308; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_310 = 10'h136 == index ? 32'h67756265 : _GEN_309; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_311 = 10'h137 == index ? 32'h3331302d : _GEN_310; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_312 = 10'h138 == index ? 32'h0 : _GEN_311; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_313 = 10'h139 == index ? 32'h3000000 : _GEN_312; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_314 = 10'h13a == index ? 32'h4000000 : _GEN_313; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_315 = 10'h13b == index ? 32'h9d010000 : _GEN_314; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_316 = 10'h13c == index ? 32'h696d64 : _GEN_315; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_317 = 10'h13d == index ? 32'h3000000 : _GEN_316; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_318 = 10'h13e == index ? 32'h8000000 : _GEN_317; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_319 = 10'h13f == index ? 32'h7f010000 : _GEN_318; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_320 = 10'h140 == index ? 32'h2000000 : _GEN_319; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_321 = 10'h141 == index ? 32'hffff0000 : _GEN_320; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_322 = 10'h142 == index ? 32'h3000000 : _GEN_321; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_323 = 10'h143 == index ? 32'h8000000 : _GEN_322; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_324 = 10'h144 == index ? 32'h7010000 : _GEN_323; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_325 = 10'h145 == index ? 32'h0 : _GEN_324; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_326 = 10'h146 == index ? 32'h100000 : _GEN_325; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_327 = 10'h147 == index ? 32'h3000000 : _GEN_326; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_328 = 10'h148 == index ? 32'h8000000 : _GEN_327; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_329 = 10'h149 == index ? 32'h93010000 : _GEN_328; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_330 = 10'h14a == index ? 32'h746e6f63 : _GEN_329; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_331 = 10'h14b == index ? 32'h6c6f72 : _GEN_330; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_332 = 10'h14c == index ? 32'h2000000 : _GEN_331; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_333 = 10'h14d == index ? 32'h1000000 : _GEN_332; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_334 = 10'h14e == index ? 32'h6f727265 : _GEN_333; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_335 = 10'h14f == index ? 32'h65642d72 : _GEN_334; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_336 = 10'h150 == index ? 32'h65636976 : _GEN_335; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_337 = 10'h151 == index ? 32'h30303340 : _GEN_336; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_338 = 10'h152 == index ? 32'h30 : _GEN_337; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_339 = 10'h153 == index ? 32'h3000000 : _GEN_338; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_340 = 10'h154 == index ? 32'he000000 : _GEN_339; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_341 = 10'h155 == index ? 32'h1b000000 : _GEN_340; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_342 = 10'h156 == index ? 32'h69666973 : _GEN_341; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_343 = 10'h157 == index ? 32'h652c6576 : _GEN_342; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_344 = 10'h158 == index ? 32'h726f7272 : _GEN_343; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_345 = 10'h159 == index ? 32'h30 : _GEN_344; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_346 = 10'h15a == index ? 32'h3000000 : _GEN_345; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_347 = 10'h15b == index ? 32'h8000000 : _GEN_346; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_348 = 10'h15c == index ? 32'h7010000 : _GEN_347; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_349 = 10'h15d == index ? 32'h300000 : _GEN_348; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_350 = 10'h15e == index ? 32'h100000 : _GEN_349; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_351 = 10'h15f == index ? 32'h2000000 : _GEN_350; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_352 = 10'h160 == index ? 32'h1000000 : _GEN_351; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_353 = 10'h161 == index ? 32'h65747865 : _GEN_352; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_354 = 10'h162 == index ? 32'h6c616e72 : _GEN_353; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_355 = 10'h163 == index ? 32'h746e692d : _GEN_354; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_356 = 10'h164 == index ? 32'h75727265 : _GEN_355; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_357 = 10'h165 == index ? 32'h737470 : _GEN_356; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_358 = 10'h166 == index ? 32'h3000000 : _GEN_357; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_359 = 10'h167 == index ? 32'h4000000 : _GEN_358; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_360 = 10'h168 == index ? 32'haa010000 : _GEN_359; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_361 = 10'h169 == index ? 32'h3000000 : _GEN_360; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_362 = 10'h16a == index ? 32'h3000000 : _GEN_361; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_363 = 10'h16b == index ? 32'h8000000 : _GEN_362; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_364 = 10'h16c == index ? 32'hbb010000 : _GEN_363; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_365 = 10'h16d == index ? 32'h1000000 : _GEN_364; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_366 = 10'h16e == index ? 32'h2000000 : _GEN_365; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_367 = 10'h16f == index ? 32'h2000000 : _GEN_366; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_368 = 10'h170 == index ? 32'h1000000 : _GEN_367; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_369 = 10'h171 == index ? 32'h65746e69 : _GEN_368; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_370 = 10'h172 == index ? 32'h70757272 : _GEN_369; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_371 = 10'h173 == index ? 32'h6f632d74 : _GEN_370; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_372 = 10'h174 == index ? 32'h6f72746e : _GEN_371; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_373 = 10'h175 == index ? 32'h72656c6c : _GEN_372; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_374 = 10'h176 == index ? 32'h30306340 : _GEN_373; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_375 = 10'h177 == index ? 32'h30303030 : _GEN_374; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_376 = 10'h178 == index ? 32'h0 : _GEN_375; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_377 = 10'h179 == index ? 32'h3000000 : _GEN_376; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_378 = 10'h17a == index ? 32'h4000000 : _GEN_377; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_379 = 10'h17b == index ? 32'h4a010000 : _GEN_378; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_380 = 10'h17c == index ? 32'h1000000 : _GEN_379; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_381 = 10'h17d == index ? 32'h3000000 : _GEN_380; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_382 = 10'h17e == index ? 32'hc000000 : _GEN_381; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_383 = 10'h17f == index ? 32'h1b000000 : _GEN_382; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_384 = 10'h180 == index ? 32'h63736972 : _GEN_383; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_385 = 10'h181 == index ? 32'h6c702c76 : _GEN_384; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_386 = 10'h182 == index ? 32'h306369 : _GEN_385; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_387 = 10'h183 == index ? 32'h3000000 : _GEN_386; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_388 = 10'h184 == index ? 32'h0 : _GEN_387; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_389 = 10'h185 == index ? 32'h5b010000 : _GEN_388; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_390 = 10'h186 == index ? 32'h3000000 : _GEN_389; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_391 = 10'h187 == index ? 32'h10000000 : _GEN_390; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_392 = 10'h188 == index ? 32'h7f010000 : _GEN_391; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_393 = 10'h189 == index ? 32'h2000000 : _GEN_392; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_394 = 10'h18a == index ? 32'hb000000 : _GEN_393; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_395 = 10'h18b == index ? 32'h2000000 : _GEN_394; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_396 = 10'h18c == index ? 32'h9000000 : _GEN_395; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_397 = 10'h18d == index ? 32'h3000000 : _GEN_396; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_398 = 10'h18e == index ? 32'h8000000 : _GEN_397; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_399 = 10'h18f == index ? 32'h7010000 : _GEN_398; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_400 = 10'h190 == index ? 32'hc : _GEN_399; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_401 = 10'h191 == index ? 32'h4 : _GEN_400; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_402 = 10'h192 == index ? 32'h3000000 : _GEN_401; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_403 = 10'h193 == index ? 32'h8000000 : _GEN_402; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_404 = 10'h194 == index ? 32'h93010000 : _GEN_403; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_405 = 10'h195 == index ? 32'h746e6f63 : _GEN_404; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_406 = 10'h196 == index ? 32'h6c6f72 : _GEN_405; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_407 = 10'h197 == index ? 32'h3000000 : _GEN_406; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_408 = 10'h198 == index ? 32'h4000000 : _GEN_407; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_409 = 10'h199 == index ? 32'hc6010000 : _GEN_408; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_410 = 10'h19a == index ? 32'h3000000 : _GEN_409; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_411 = 10'h19b == index ? 32'h3000000 : _GEN_410; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_412 = 10'h19c == index ? 32'h4000000 : _GEN_411; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_413 = 10'h19d == index ? 32'hd9010000 : _GEN_412; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_414 = 10'h19e == index ? 32'h2000000 : _GEN_413; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_415 = 10'h19f == index ? 32'h3000000 : _GEN_414; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_416 = 10'h1a0 == index ? 32'h4000000 : _GEN_415; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_417 = 10'h1a1 == index ? 32'h70010000 : _GEN_416; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_418 = 10'h1a2 == index ? 32'h3000000 : _GEN_417; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_419 = 10'h1a3 == index ? 32'h2000000 : _GEN_418; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_420 = 10'h1a4 == index ? 32'h1000000 : _GEN_419; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_421 = 10'h1a5 == index ? 32'h6f696d6d : _GEN_420; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_422 = 10'h1a6 == index ? 32'h726f702d : _GEN_421; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_423 = 10'h1a7 == index ? 32'h78612d74 : _GEN_422; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_424 = 10'h1a8 == index ? 32'h36403469 : _GEN_423; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_425 = 10'h1a9 == index ? 32'h30303030 : _GEN_424; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_426 = 10'h1aa == index ? 32'h303030 : _GEN_425; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_427 = 10'h1ab == index ? 32'h3000000 : _GEN_426; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_428 = 10'h1ac == index ? 32'h4000000 : _GEN_427; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_429 = 10'h1ad == index ? 32'h0 : _GEN_428; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_430 = 10'h1ae == index ? 32'h1000000 : _GEN_429; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_431 = 10'h1af == index ? 32'h3000000 : _GEN_430; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_432 = 10'h1b0 == index ? 32'h4000000 : _GEN_431; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_433 = 10'h1b1 == index ? 32'hf000000 : _GEN_432; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_434 = 10'h1b2 == index ? 32'h1000000 : _GEN_433; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_435 = 10'h1b3 == index ? 32'h3000000 : _GEN_434; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_436 = 10'h1b4 == index ? 32'hb000000 : _GEN_435; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_437 = 10'h1b5 == index ? 32'h1b000000 : _GEN_436; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_438 = 10'h1b6 == index ? 32'h706d6973 : _GEN_437; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_439 = 10'h1b7 == index ? 32'h622d656c : _GEN_438; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_440 = 10'h1b8 == index ? 32'h7375 : _GEN_439; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_441 = 10'h1b9 == index ? 32'h3000000 : _GEN_440; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_442 = 10'h1ba == index ? 32'hc000000 : _GEN_441; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_443 = 10'h1bb == index ? 32'h78010000 : _GEN_442; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_444 = 10'h1bc == index ? 32'h60 : _GEN_443; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_445 = 10'h1bd == index ? 32'h60 : _GEN_444; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_446 = 10'h1be == index ? 32'h20 : _GEN_445; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_447 = 10'h1bf == index ? 32'h2000000 : _GEN_446; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_448 = 10'h1c0 == index ? 32'h1000000 : _GEN_447; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_449 = 10'h1c1 == index ? 32'h406d6f72 : _GEN_448; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_450 = 10'h1c2 == index ? 32'h30303031 : _GEN_449; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_451 = 10'h1c3 == index ? 32'h30 : _GEN_450; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_452 = 10'h1c4 == index ? 32'h3000000 : _GEN_451; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_453 = 10'h1c5 == index ? 32'hc000000 : _GEN_452; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_454 = 10'h1c6 == index ? 32'h1b000000 : _GEN_453; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_455 = 10'h1c7 == index ? 32'h69666973 : _GEN_454; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_456 = 10'h1c8 == index ? 32'h722c6576 : _GEN_455; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_457 = 10'h1c9 == index ? 32'h306d6f : _GEN_456; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_458 = 10'h1ca == index ? 32'h3000000 : _GEN_457; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_459 = 10'h1cb == index ? 32'h8000000 : _GEN_458; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_460 = 10'h1cc == index ? 32'h7010000 : _GEN_459; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_461 = 10'h1cd == index ? 32'h100 : _GEN_460; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_462 = 10'h1ce == index ? 32'h100 : _GEN_461; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_463 = 10'h1cf == index ? 32'h3000000 : _GEN_462; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_464 = 10'h1d0 == index ? 32'h4000000 : _GEN_463; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_465 = 10'h1d1 == index ? 32'h93010000 : _GEN_464; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_466 = 10'h1d2 == index ? 32'h6d656d : _GEN_465; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_467 = 10'h1d3 == index ? 32'h2000000 : _GEN_466; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_468 = 10'h1d4 == index ? 32'h2000000 : _GEN_467; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_469 = 10'h1d5 == index ? 32'h2000000 : _GEN_468; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_470 = 10'h1d6 == index ? 32'h9000000 : _GEN_469; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_471 = 10'h1d7 == index ? 32'h64646123 : _GEN_470; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_472 = 10'h1d8 == index ? 32'h73736572 : _GEN_471; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_473 = 10'h1d9 == index ? 32'h6c65632d : _GEN_472; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_474 = 10'h1da == index ? 32'h2300736c : _GEN_473; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_475 = 10'h1db == index ? 32'h657a6973 : _GEN_474; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_476 = 10'h1dc == index ? 32'h6c65632d : _GEN_475; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_477 = 10'h1dd == index ? 32'h6300736c : _GEN_476; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_478 = 10'h1de == index ? 32'h61706d6f : _GEN_477; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_479 = 10'h1df == index ? 32'h6c626974 : _GEN_478; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_480 = 10'h1e0 == index ? 32'h6f6d0065 : _GEN_479; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_481 = 10'h1e1 == index ? 32'h6c6564 : _GEN_480; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_482 = 10'h1e2 == index ? 32'h636f6c63 : _GEN_481; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_483 = 10'h1e3 == index ? 32'h72662d6b : _GEN_482; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_484 = 10'h1e4 == index ? 32'h65757165 : _GEN_483; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_485 = 10'h1e5 == index ? 32'h79636e : _GEN_484; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_486 = 10'h1e6 == index ? 32'h61632d64 : _GEN_485; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_487 = 10'h1e7 == index ? 32'h2d656863 : _GEN_486; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_488 = 10'h1e8 == index ? 32'h636f6c62 : _GEN_487; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_489 = 10'h1e9 == index ? 32'h69732d6b : _GEN_488; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_490 = 10'h1ea == index ? 32'h6400657a : _GEN_489; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_491 = 10'h1eb == index ? 32'h6361632d : _GEN_490; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_492 = 10'h1ec == index ? 32'h732d6568 : _GEN_491; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_493 = 10'h1ed == index ? 32'h737465 : _GEN_492; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_494 = 10'h1ee == index ? 32'h61632d64 : _GEN_493; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_495 = 10'h1ef == index ? 32'h2d656863 : _GEN_494; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_496 = 10'h1f0 == index ? 32'h657a6973 : _GEN_495; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_497 = 10'h1f1 == index ? 32'h742d6400 : _GEN_496; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_498 = 10'h1f2 == index ? 32'h732d626c : _GEN_497; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_499 = 10'h1f3 == index ? 32'h737465 : _GEN_498; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_500 = 10'h1f4 == index ? 32'h6c742d64 : _GEN_499; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_501 = 10'h1f5 == index ? 32'h69732d62 : _GEN_500; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_502 = 10'h1f6 == index ? 32'h6400657a : _GEN_501; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_503 = 10'h1f7 == index ? 32'h63697665 : _GEN_502; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_504 = 10'h1f8 == index ? 32'h79745f65 : _GEN_503; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_505 = 10'h1f9 == index ? 32'h68006570 : _GEN_504; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_506 = 10'h1fa == index ? 32'h77647261 : _GEN_505; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_507 = 10'h1fb == index ? 32'h2d657261 : _GEN_506; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_508 = 10'h1fc == index ? 32'h63657865 : _GEN_507; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_509 = 10'h1fd == index ? 32'h6572622d : _GEN_508; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_510 = 10'h1fe == index ? 32'h6f706b61 : _GEN_509; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_511 = 10'h1ff == index ? 32'h2d746e69 : _GEN_510; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_512 = 10'h200 == index ? 32'h6e756f63 : _GEN_511; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_513 = 10'h201 == index ? 32'h2d690074 : _GEN_512; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_514 = 10'h202 == index ? 32'h68636163 : _GEN_513; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_515 = 10'h203 == index ? 32'h6c622d65 : _GEN_514; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_516 = 10'h204 == index ? 32'h2d6b636f : _GEN_515; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_517 = 10'h205 == index ? 32'h657a6973 : _GEN_516; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_518 = 10'h206 == index ? 32'h632d6900 : _GEN_517; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_519 = 10'h207 == index ? 32'h65686361 : _GEN_518; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_520 = 10'h208 == index ? 32'h7465732d : _GEN_519; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_521 = 10'h209 == index ? 32'h2d690073 : _GEN_520; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_522 = 10'h20a == index ? 32'h68636163 : _GEN_521; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_523 = 10'h20b == index ? 32'h69732d65 : _GEN_522; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_524 = 10'h20c == index ? 32'h6900657a : _GEN_523; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_525 = 10'h20d == index ? 32'h626c742d : _GEN_524; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_526 = 10'h20e == index ? 32'h7465732d : _GEN_525; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_527 = 10'h20f == index ? 32'h2d690073 : _GEN_526; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_528 = 10'h210 == index ? 32'h2d626c74 : _GEN_527; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_529 = 10'h211 == index ? 32'h657a6973 : _GEN_528; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_530 = 10'h212 == index ? 32'h756d6d00 : _GEN_529; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_531 = 10'h213 == index ? 32'h7079742d : _GEN_530; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_532 = 10'h214 == index ? 32'h656e0065 : _GEN_531; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_533 = 10'h215 == index ? 32'h6c2d7478 : _GEN_532; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_534 = 10'h216 == index ? 32'h6c657665 : _GEN_533; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_535 = 10'h217 == index ? 32'h6361632d : _GEN_534; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_536 = 10'h218 == index ? 32'h72006568 : _GEN_535; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_537 = 10'h219 == index ? 32'h72006765 : _GEN_536; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_538 = 10'h21a == index ? 32'h76637369 : _GEN_537; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_539 = 10'h21b == index ? 32'h6173692c : _GEN_538; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_540 = 10'h21c == index ? 32'h73697200 : _GEN_539; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_541 = 10'h21d == index ? 32'h702c7663 : _GEN_540; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_542 = 10'h21e == index ? 32'h6572706d : _GEN_541; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_543 = 10'h21f == index ? 32'h6e6f6967 : _GEN_542; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_544 = 10'h220 == index ? 32'h74730073 : _GEN_543; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_545 = 10'h221 == index ? 32'h73757461 : _GEN_544; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_546 = 10'h222 == index ? 32'h6d697400 : _GEN_545; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_547 = 10'h223 == index ? 32'h73616265 : _GEN_546; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_548 = 10'h224 == index ? 32'h72662d65 : _GEN_547; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_549 = 10'h225 == index ? 32'h65757165 : _GEN_548; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_550 = 10'h226 == index ? 32'h79636e : _GEN_549; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_551 = 10'h227 == index ? 32'h2d626c74 : _GEN_550; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_552 = 10'h228 == index ? 32'h696c7073 : _GEN_551; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_553 = 10'h229 == index ? 32'h69230074 : _GEN_552; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_554 = 10'h22a == index ? 32'h7265746e : _GEN_553; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_555 = 10'h22b == index ? 32'h74707572 : _GEN_554; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_556 = 10'h22c == index ? 32'h6c65632d : _GEN_555; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_557 = 10'h22d == index ? 32'h6900736c : _GEN_556; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_558 = 10'h22e == index ? 32'h7265746e : _GEN_557; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_559 = 10'h22f == index ? 32'h74707572 : _GEN_558; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_560 = 10'h230 == index ? 32'h6e6f632d : _GEN_559; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_561 = 10'h231 == index ? 32'h6c6f7274 : _GEN_560; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_562 = 10'h232 == index ? 32'h72656c : _GEN_561; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_563 = 10'h233 == index ? 32'h6e616870 : _GEN_562; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_564 = 10'h234 == index ? 32'h656c64 : _GEN_563; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_565 = 10'h235 == index ? 32'h676e6172 : _GEN_564; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_566 = 10'h236 == index ? 32'h69007365 : _GEN_565; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_567 = 10'h237 == index ? 32'h7265746e : _GEN_566; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_568 = 10'h238 == index ? 32'h74707572 : _GEN_567; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_569 = 10'h239 == index ? 32'h78652d73 : _GEN_568; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_570 = 10'h23a == index ? 32'h646e6574 : _GEN_569; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_571 = 10'h23b == index ? 32'h72006465 : _GEN_570; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_572 = 10'h23c == index ? 32'h6e2d6765 : _GEN_571; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_573 = 10'h23d == index ? 32'h73656d61 : _GEN_572; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_574 = 10'h23e == index ? 32'h62656400 : _GEN_573; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_575 = 10'h23f == index ? 32'h612d6775 : _GEN_574; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_576 = 10'h240 == index ? 32'h63617474 : _GEN_575; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_577 = 10'h241 == index ? 32'h6e690068 : _GEN_576; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_578 = 10'h242 == index ? 32'h72726574 : _GEN_577; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_579 = 10'h243 == index ? 32'h2d747075 : _GEN_578; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_580 = 10'h244 == index ? 32'h65726170 : _GEN_579; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_581 = 10'h245 == index ? 32'h6900746e : _GEN_580; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_582 = 10'h246 == index ? 32'h7265746e : _GEN_581; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_583 = 10'h247 == index ? 32'h74707572 : _GEN_582; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_584 = 10'h248 == index ? 32'h69720073 : _GEN_583; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_585 = 10'h249 == index ? 32'h2c766373 : _GEN_584; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_586 = 10'h24a == index ? 32'h2d78616d : _GEN_585; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_587 = 10'h24b == index ? 32'h6f697270 : _GEN_586; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_588 = 10'h24c == index ? 32'h79746972 : _GEN_587; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_589 = 10'h24d == index ? 32'h73697200 : _GEN_588; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_590 = 10'h24e == index ? 32'h6e2c7663 : _GEN_589; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_591 = 10'h24f == index ? 32'h766564 : _GEN_590; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_592 = 10'h250 == index ? 32'h0 : _GEN_591; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_593 = 10'h251 == index ? 32'h0 : _GEN_592; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_594 = 10'h252 == index ? 32'h0 : _GEN_593; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_595 = 10'h253 == index ? 32'h0 : _GEN_594; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_596 = 10'h254 == index ? 32'h0 : _GEN_595; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_597 = 10'h255 == index ? 32'h0 : _GEN_596; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_598 = 10'h256 == index ? 32'h0 : _GEN_597; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_599 = 10'h257 == index ? 32'h0 : _GEN_598; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_600 = 10'h258 == index ? 32'h0 : _GEN_599; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_601 = 10'h259 == index ? 32'h0 : _GEN_600; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_602 = 10'h25a == index ? 32'h0 : _GEN_601; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_603 = 10'h25b == index ? 32'h0 : _GEN_602; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_604 = 10'h25c == index ? 32'h0 : _GEN_603; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_605 = 10'h25d == index ? 32'h0 : _GEN_604; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_606 = 10'h25e == index ? 32'h0 : _GEN_605; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_607 = 10'h25f == index ? 32'h0 : _GEN_606; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_608 = 10'h260 == index ? 32'h0 : _GEN_607; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_609 = 10'h261 == index ? 32'h0 : _GEN_608; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_610 = 10'h262 == index ? 32'h0 : _GEN_609; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_611 = 10'h263 == index ? 32'h0 : _GEN_610; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_612 = 10'h264 == index ? 32'h0 : _GEN_611; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_613 = 10'h265 == index ? 32'h0 : _GEN_612; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_614 = 10'h266 == index ? 32'h0 : _GEN_613; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_615 = 10'h267 == index ? 32'h0 : _GEN_614; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_616 = 10'h268 == index ? 32'h0 : _GEN_615; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_617 = 10'h269 == index ? 32'h0 : _GEN_616; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_618 = 10'h26a == index ? 32'h0 : _GEN_617; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_619 = 10'h26b == index ? 32'h0 : _GEN_618; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_620 = 10'h26c == index ? 32'h0 : _GEN_619; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_621 = 10'h26d == index ? 32'h0 : _GEN_620; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_622 = 10'h26e == index ? 32'h0 : _GEN_621; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_623 = 10'h26f == index ? 32'h0 : _GEN_622; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_624 = 10'h270 == index ? 32'h0 : _GEN_623; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_625 = 10'h271 == index ? 32'h0 : _GEN_624; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_626 = 10'h272 == index ? 32'h0 : _GEN_625; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_627 = 10'h273 == index ? 32'h0 : _GEN_626; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_628 = 10'h274 == index ? 32'h0 : _GEN_627; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_629 = 10'h275 == index ? 32'h0 : _GEN_628; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_630 = 10'h276 == index ? 32'h0 : _GEN_629; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_631 = 10'h277 == index ? 32'h0 : _GEN_630; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_632 = 10'h278 == index ? 32'h0 : _GEN_631; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_633 = 10'h279 == index ? 32'h0 : _GEN_632; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_634 = 10'h27a == index ? 32'h0 : _GEN_633; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_635 = 10'h27b == index ? 32'h0 : _GEN_634; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_636 = 10'h27c == index ? 32'h0 : _GEN_635; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_637 = 10'h27d == index ? 32'h0 : _GEN_636; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_638 = 10'h27e == index ? 32'h0 : _GEN_637; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_639 = 10'h27f == index ? 32'h0 : _GEN_638; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_640 = 10'h280 == index ? 32'h0 : _GEN_639; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_641 = 10'h281 == index ? 32'h0 : _GEN_640; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_642 = 10'h282 == index ? 32'h0 : _GEN_641; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_643 = 10'h283 == index ? 32'h0 : _GEN_642; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_644 = 10'h284 == index ? 32'h0 : _GEN_643; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_645 = 10'h285 == index ? 32'h0 : _GEN_644; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_646 = 10'h286 == index ? 32'h0 : _GEN_645; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_647 = 10'h287 == index ? 32'h0 : _GEN_646; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_648 = 10'h288 == index ? 32'h0 : _GEN_647; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_649 = 10'h289 == index ? 32'h0 : _GEN_648; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_650 = 10'h28a == index ? 32'h0 : _GEN_649; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_651 = 10'h28b == index ? 32'h0 : _GEN_650; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_652 = 10'h28c == index ? 32'h0 : _GEN_651; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_653 = 10'h28d == index ? 32'h0 : _GEN_652; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_654 = 10'h28e == index ? 32'h0 : _GEN_653; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_655 = 10'h28f == index ? 32'h0 : _GEN_654; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_656 = 10'h290 == index ? 32'h0 : _GEN_655; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_657 = 10'h291 == index ? 32'h0 : _GEN_656; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_658 = 10'h292 == index ? 32'h0 : _GEN_657; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_659 = 10'h293 == index ? 32'h0 : _GEN_658; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_660 = 10'h294 == index ? 32'h0 : _GEN_659; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_661 = 10'h295 == index ? 32'h0 : _GEN_660; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_662 = 10'h296 == index ? 32'h0 : _GEN_661; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_663 = 10'h297 == index ? 32'h0 : _GEN_662; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_664 = 10'h298 == index ? 32'h0 : _GEN_663; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_665 = 10'h299 == index ? 32'h0 : _GEN_664; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_666 = 10'h29a == index ? 32'h0 : _GEN_665; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_667 = 10'h29b == index ? 32'h0 : _GEN_666; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_668 = 10'h29c == index ? 32'h0 : _GEN_667; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_669 = 10'h29d == index ? 32'h0 : _GEN_668; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_670 = 10'h29e == index ? 32'h0 : _GEN_669; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_671 = 10'h29f == index ? 32'h0 : _GEN_670; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_672 = 10'h2a0 == index ? 32'h0 : _GEN_671; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_673 = 10'h2a1 == index ? 32'h0 : _GEN_672; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_674 = 10'h2a2 == index ? 32'h0 : _GEN_673; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_675 = 10'h2a3 == index ? 32'h0 : _GEN_674; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_676 = 10'h2a4 == index ? 32'h0 : _GEN_675; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_677 = 10'h2a5 == index ? 32'h0 : _GEN_676; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_678 = 10'h2a6 == index ? 32'h0 : _GEN_677; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_679 = 10'h2a7 == index ? 32'h0 : _GEN_678; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_680 = 10'h2a8 == index ? 32'h0 : _GEN_679; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_681 = 10'h2a9 == index ? 32'h0 : _GEN_680; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_682 = 10'h2aa == index ? 32'h0 : _GEN_681; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_683 = 10'h2ab == index ? 32'h0 : _GEN_682; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_684 = 10'h2ac == index ? 32'h0 : _GEN_683; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_685 = 10'h2ad == index ? 32'h0 : _GEN_684; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_686 = 10'h2ae == index ? 32'h0 : _GEN_685; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_687 = 10'h2af == index ? 32'h0 : _GEN_686; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_688 = 10'h2b0 == index ? 32'h0 : _GEN_687; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_689 = 10'h2b1 == index ? 32'h0 : _GEN_688; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_690 = 10'h2b2 == index ? 32'h0 : _GEN_689; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_691 = 10'h2b3 == index ? 32'h0 : _GEN_690; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_692 = 10'h2b4 == index ? 32'h0 : _GEN_691; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_693 = 10'h2b5 == index ? 32'h0 : _GEN_692; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_694 = 10'h2b6 == index ? 32'h0 : _GEN_693; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_695 = 10'h2b7 == index ? 32'h0 : _GEN_694; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_696 = 10'h2b8 == index ? 32'h0 : _GEN_695; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_697 = 10'h2b9 == index ? 32'h0 : _GEN_696; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_698 = 10'h2ba == index ? 32'h0 : _GEN_697; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_699 = 10'h2bb == index ? 32'h0 : _GEN_698; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_700 = 10'h2bc == index ? 32'h0 : _GEN_699; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_701 = 10'h2bd == index ? 32'h0 : _GEN_700; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_702 = 10'h2be == index ? 32'h0 : _GEN_701; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_703 = 10'h2bf == index ? 32'h0 : _GEN_702; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_704 = 10'h2c0 == index ? 32'h0 : _GEN_703; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_705 = 10'h2c1 == index ? 32'h0 : _GEN_704; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_706 = 10'h2c2 == index ? 32'h0 : _GEN_705; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_707 = 10'h2c3 == index ? 32'h0 : _GEN_706; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_708 = 10'h2c4 == index ? 32'h0 : _GEN_707; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_709 = 10'h2c5 == index ? 32'h0 : _GEN_708; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_710 = 10'h2c6 == index ? 32'h0 : _GEN_709; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_711 = 10'h2c7 == index ? 32'h0 : _GEN_710; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_712 = 10'h2c8 == index ? 32'h0 : _GEN_711; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_713 = 10'h2c9 == index ? 32'h0 : _GEN_712; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_714 = 10'h2ca == index ? 32'h0 : _GEN_713; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_715 = 10'h2cb == index ? 32'h0 : _GEN_714; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_716 = 10'h2cc == index ? 32'h0 : _GEN_715; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_717 = 10'h2cd == index ? 32'h0 : _GEN_716; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_718 = 10'h2ce == index ? 32'h0 : _GEN_717; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_719 = 10'h2cf == index ? 32'h0 : _GEN_718; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_720 = 10'h2d0 == index ? 32'h0 : _GEN_719; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_721 = 10'h2d1 == index ? 32'h0 : _GEN_720; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_722 = 10'h2d2 == index ? 32'h0 : _GEN_721; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_723 = 10'h2d3 == index ? 32'h0 : _GEN_722; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_724 = 10'h2d4 == index ? 32'h0 : _GEN_723; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_725 = 10'h2d5 == index ? 32'h0 : _GEN_724; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_726 = 10'h2d6 == index ? 32'h0 : _GEN_725; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_727 = 10'h2d7 == index ? 32'h0 : _GEN_726; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_728 = 10'h2d8 == index ? 32'h0 : _GEN_727; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_729 = 10'h2d9 == index ? 32'h0 : _GEN_728; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_730 = 10'h2da == index ? 32'h0 : _GEN_729; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_731 = 10'h2db == index ? 32'h0 : _GEN_730; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_732 = 10'h2dc == index ? 32'h0 : _GEN_731; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_733 = 10'h2dd == index ? 32'h0 : _GEN_732; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_734 = 10'h2de == index ? 32'h0 : _GEN_733; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_735 = 10'h2df == index ? 32'h0 : _GEN_734; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_736 = 10'h2e0 == index ? 32'h0 : _GEN_735; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_737 = 10'h2e1 == index ? 32'h0 : _GEN_736; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_738 = 10'h2e2 == index ? 32'h0 : _GEN_737; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_739 = 10'h2e3 == index ? 32'h0 : _GEN_738; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_740 = 10'h2e4 == index ? 32'h0 : _GEN_739; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_741 = 10'h2e5 == index ? 32'h0 : _GEN_740; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_742 = 10'h2e6 == index ? 32'h0 : _GEN_741; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_743 = 10'h2e7 == index ? 32'h0 : _GEN_742; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_744 = 10'h2e8 == index ? 32'h0 : _GEN_743; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_745 = 10'h2e9 == index ? 32'h0 : _GEN_744; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_746 = 10'h2ea == index ? 32'h0 : _GEN_745; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_747 = 10'h2eb == index ? 32'h0 : _GEN_746; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_748 = 10'h2ec == index ? 32'h0 : _GEN_747; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_749 = 10'h2ed == index ? 32'h0 : _GEN_748; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_750 = 10'h2ee == index ? 32'h0 : _GEN_749; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_751 = 10'h2ef == index ? 32'h0 : _GEN_750; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_752 = 10'h2f0 == index ? 32'h0 : _GEN_751; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_753 = 10'h2f1 == index ? 32'h0 : _GEN_752; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_754 = 10'h2f2 == index ? 32'h0 : _GEN_753; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_755 = 10'h2f3 == index ? 32'h0 : _GEN_754; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_756 = 10'h2f4 == index ? 32'h0 : _GEN_755; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_757 = 10'h2f5 == index ? 32'h0 : _GEN_756; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_758 = 10'h2f6 == index ? 32'h0 : _GEN_757; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_759 = 10'h2f7 == index ? 32'h0 : _GEN_758; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_760 = 10'h2f8 == index ? 32'h0 : _GEN_759; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_761 = 10'h2f9 == index ? 32'h0 : _GEN_760; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_762 = 10'h2fa == index ? 32'h0 : _GEN_761; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_763 = 10'h2fb == index ? 32'h0 : _GEN_762; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_764 = 10'h2fc == index ? 32'h0 : _GEN_763; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_765 = 10'h2fd == index ? 32'h0 : _GEN_764; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_766 = 10'h2fe == index ? 32'h0 : _GEN_765; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_767 = 10'h2ff == index ? 32'h0 : _GEN_766; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_768 = 10'h300 == index ? 32'h0 : _GEN_767; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_769 = 10'h301 == index ? 32'h0 : _GEN_768; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_770 = 10'h302 == index ? 32'h0 : _GEN_769; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_771 = 10'h303 == index ? 32'h0 : _GEN_770; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_772 = 10'h304 == index ? 32'h0 : _GEN_771; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_773 = 10'h305 == index ? 32'h0 : _GEN_772; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_774 = 10'h306 == index ? 32'h0 : _GEN_773; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_775 = 10'h307 == index ? 32'h0 : _GEN_774; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_776 = 10'h308 == index ? 32'h0 : _GEN_775; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_777 = 10'h309 == index ? 32'h0 : _GEN_776; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_778 = 10'h30a == index ? 32'h0 : _GEN_777; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_779 = 10'h30b == index ? 32'h0 : _GEN_778; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_780 = 10'h30c == index ? 32'h0 : _GEN_779; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_781 = 10'h30d == index ? 32'h0 : _GEN_780; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_782 = 10'h30e == index ? 32'h0 : _GEN_781; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_783 = 10'h30f == index ? 32'h0 : _GEN_782; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_784 = 10'h310 == index ? 32'h0 : _GEN_783; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_785 = 10'h311 == index ? 32'h0 : _GEN_784; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_786 = 10'h312 == index ? 32'h0 : _GEN_785; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_787 = 10'h313 == index ? 32'h0 : _GEN_786; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_788 = 10'h314 == index ? 32'h0 : _GEN_787; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_789 = 10'h315 == index ? 32'h0 : _GEN_788; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_790 = 10'h316 == index ? 32'h0 : _GEN_789; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_791 = 10'h317 == index ? 32'h0 : _GEN_790; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_792 = 10'h318 == index ? 32'h0 : _GEN_791; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_793 = 10'h319 == index ? 32'h0 : _GEN_792; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_794 = 10'h31a == index ? 32'h0 : _GEN_793; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_795 = 10'h31b == index ? 32'h0 : _GEN_794; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_796 = 10'h31c == index ? 32'h0 : _GEN_795; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_797 = 10'h31d == index ? 32'h0 : _GEN_796; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_798 = 10'h31e == index ? 32'h0 : _GEN_797; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_799 = 10'h31f == index ? 32'h0 : _GEN_798; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_800 = 10'h320 == index ? 32'h0 : _GEN_799; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_801 = 10'h321 == index ? 32'h0 : _GEN_800; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_802 = 10'h322 == index ? 32'h0 : _GEN_801; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_803 = 10'h323 == index ? 32'h0 : _GEN_802; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_804 = 10'h324 == index ? 32'h0 : _GEN_803; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_805 = 10'h325 == index ? 32'h0 : _GEN_804; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_806 = 10'h326 == index ? 32'h0 : _GEN_805; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_807 = 10'h327 == index ? 32'h0 : _GEN_806; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_808 = 10'h328 == index ? 32'h0 : _GEN_807; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_809 = 10'h329 == index ? 32'h0 : _GEN_808; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_810 = 10'h32a == index ? 32'h0 : _GEN_809; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_811 = 10'h32b == index ? 32'h0 : _GEN_810; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_812 = 10'h32c == index ? 32'h0 : _GEN_811; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_813 = 10'h32d == index ? 32'h0 : _GEN_812; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_814 = 10'h32e == index ? 32'h0 : _GEN_813; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_815 = 10'h32f == index ? 32'h0 : _GEN_814; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_816 = 10'h330 == index ? 32'h0 : _GEN_815; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_817 = 10'h331 == index ? 32'h0 : _GEN_816; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_818 = 10'h332 == index ? 32'h0 : _GEN_817; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_819 = 10'h333 == index ? 32'h0 : _GEN_818; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_820 = 10'h334 == index ? 32'h0 : _GEN_819; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_821 = 10'h335 == index ? 32'h0 : _GEN_820; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_822 = 10'h336 == index ? 32'h0 : _GEN_821; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_823 = 10'h337 == index ? 32'h0 : _GEN_822; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_824 = 10'h338 == index ? 32'h0 : _GEN_823; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_825 = 10'h339 == index ? 32'h0 : _GEN_824; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_826 = 10'h33a == index ? 32'h0 : _GEN_825; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_827 = 10'h33b == index ? 32'h0 : _GEN_826; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_828 = 10'h33c == index ? 32'h0 : _GEN_827; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_829 = 10'h33d == index ? 32'h0 : _GEN_828; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_830 = 10'h33e == index ? 32'h0 : _GEN_829; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_831 = 10'h33f == index ? 32'h0 : _GEN_830; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_832 = 10'h340 == index ? 32'h0 : _GEN_831; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_833 = 10'h341 == index ? 32'h0 : _GEN_832; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_834 = 10'h342 == index ? 32'h0 : _GEN_833; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_835 = 10'h343 == index ? 32'h0 : _GEN_834; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_836 = 10'h344 == index ? 32'h0 : _GEN_835; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_837 = 10'h345 == index ? 32'h0 : _GEN_836; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_838 = 10'h346 == index ? 32'h0 : _GEN_837; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_839 = 10'h347 == index ? 32'h0 : _GEN_838; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_840 = 10'h348 == index ? 32'h0 : _GEN_839; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_841 = 10'h349 == index ? 32'h0 : _GEN_840; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_842 = 10'h34a == index ? 32'h0 : _GEN_841; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_843 = 10'h34b == index ? 32'h0 : _GEN_842; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_844 = 10'h34c == index ? 32'h0 : _GEN_843; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_845 = 10'h34d == index ? 32'h0 : _GEN_844; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_846 = 10'h34e == index ? 32'h0 : _GEN_845; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_847 = 10'h34f == index ? 32'h0 : _GEN_846; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_848 = 10'h350 == index ? 32'h0 : _GEN_847; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_849 = 10'h351 == index ? 32'h0 : _GEN_848; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_850 = 10'h352 == index ? 32'h0 : _GEN_849; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_851 = 10'h353 == index ? 32'h0 : _GEN_850; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_852 = 10'h354 == index ? 32'h0 : _GEN_851; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_853 = 10'h355 == index ? 32'h0 : _GEN_852; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_854 = 10'h356 == index ? 32'h0 : _GEN_853; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_855 = 10'h357 == index ? 32'h0 : _GEN_854; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_856 = 10'h358 == index ? 32'h0 : _GEN_855; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_857 = 10'h359 == index ? 32'h0 : _GEN_856; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_858 = 10'h35a == index ? 32'h0 : _GEN_857; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_859 = 10'h35b == index ? 32'h0 : _GEN_858; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_860 = 10'h35c == index ? 32'h0 : _GEN_859; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_861 = 10'h35d == index ? 32'h0 : _GEN_860; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_862 = 10'h35e == index ? 32'h0 : _GEN_861; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_863 = 10'h35f == index ? 32'h0 : _GEN_862; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_864 = 10'h360 == index ? 32'h0 : _GEN_863; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_865 = 10'h361 == index ? 32'h0 : _GEN_864; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_866 = 10'h362 == index ? 32'h0 : _GEN_865; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_867 = 10'h363 == index ? 32'h0 : _GEN_866; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_868 = 10'h364 == index ? 32'h0 : _GEN_867; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_869 = 10'h365 == index ? 32'h0 : _GEN_868; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_870 = 10'h366 == index ? 32'h0 : _GEN_869; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_871 = 10'h367 == index ? 32'h0 : _GEN_870; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_872 = 10'h368 == index ? 32'h0 : _GEN_871; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_873 = 10'h369 == index ? 32'h0 : _GEN_872; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_874 = 10'h36a == index ? 32'h0 : _GEN_873; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_875 = 10'h36b == index ? 32'h0 : _GEN_874; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_876 = 10'h36c == index ? 32'h0 : _GEN_875; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_877 = 10'h36d == index ? 32'h0 : _GEN_876; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_878 = 10'h36e == index ? 32'h0 : _GEN_877; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_879 = 10'h36f == index ? 32'h0 : _GEN_878; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_880 = 10'h370 == index ? 32'h0 : _GEN_879; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_881 = 10'h371 == index ? 32'h0 : _GEN_880; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_882 = 10'h372 == index ? 32'h0 : _GEN_881; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_883 = 10'h373 == index ? 32'h0 : _GEN_882; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_884 = 10'h374 == index ? 32'h0 : _GEN_883; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_885 = 10'h375 == index ? 32'h0 : _GEN_884; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_886 = 10'h376 == index ? 32'h0 : _GEN_885; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_887 = 10'h377 == index ? 32'h0 : _GEN_886; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_888 = 10'h378 == index ? 32'h0 : _GEN_887; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_889 = 10'h379 == index ? 32'h0 : _GEN_888; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_890 = 10'h37a == index ? 32'h0 : _GEN_889; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_891 = 10'h37b == index ? 32'h0 : _GEN_890; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_892 = 10'h37c == index ? 32'h0 : _GEN_891; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_893 = 10'h37d == index ? 32'h0 : _GEN_892; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_894 = 10'h37e == index ? 32'h0 : _GEN_893; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_895 = 10'h37f == index ? 32'h0 : _GEN_894; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_896 = 10'h380 == index ? 32'h0 : _GEN_895; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_897 = 10'h381 == index ? 32'h0 : _GEN_896; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_898 = 10'h382 == index ? 32'h0 : _GEN_897; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_899 = 10'h383 == index ? 32'h0 : _GEN_898; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_900 = 10'h384 == index ? 32'h0 : _GEN_899; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_901 = 10'h385 == index ? 32'h0 : _GEN_900; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_902 = 10'h386 == index ? 32'h0 : _GEN_901; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_903 = 10'h387 == index ? 32'h0 : _GEN_902; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_904 = 10'h388 == index ? 32'h0 : _GEN_903; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_905 = 10'h389 == index ? 32'h0 : _GEN_904; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_906 = 10'h38a == index ? 32'h0 : _GEN_905; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_907 = 10'h38b == index ? 32'h0 : _GEN_906; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_908 = 10'h38c == index ? 32'h0 : _GEN_907; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_909 = 10'h38d == index ? 32'h0 : _GEN_908; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_910 = 10'h38e == index ? 32'h0 : _GEN_909; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_911 = 10'h38f == index ? 32'h0 : _GEN_910; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_912 = 10'h390 == index ? 32'h0 : _GEN_911; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_913 = 10'h391 == index ? 32'h0 : _GEN_912; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_914 = 10'h392 == index ? 32'h0 : _GEN_913; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_915 = 10'h393 == index ? 32'h0 : _GEN_914; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_916 = 10'h394 == index ? 32'h0 : _GEN_915; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_917 = 10'h395 == index ? 32'h0 : _GEN_916; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_918 = 10'h396 == index ? 32'h0 : _GEN_917; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_919 = 10'h397 == index ? 32'h0 : _GEN_918; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_920 = 10'h398 == index ? 32'h0 : _GEN_919; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_921 = 10'h399 == index ? 32'h0 : _GEN_920; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_922 = 10'h39a == index ? 32'h0 : _GEN_921; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_923 = 10'h39b == index ? 32'h0 : _GEN_922; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_924 = 10'h39c == index ? 32'h0 : _GEN_923; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_925 = 10'h39d == index ? 32'h0 : _GEN_924; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_926 = 10'h39e == index ? 32'h0 : _GEN_925; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_927 = 10'h39f == index ? 32'h0 : _GEN_926; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_928 = 10'h3a0 == index ? 32'h0 : _GEN_927; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_929 = 10'h3a1 == index ? 32'h0 : _GEN_928; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_930 = 10'h3a2 == index ? 32'h0 : _GEN_929; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_931 = 10'h3a3 == index ? 32'h0 : _GEN_930; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_932 = 10'h3a4 == index ? 32'h0 : _GEN_931; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_933 = 10'h3a5 == index ? 32'h0 : _GEN_932; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_934 = 10'h3a6 == index ? 32'h0 : _GEN_933; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_935 = 10'h3a7 == index ? 32'h0 : _GEN_934; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_936 = 10'h3a8 == index ? 32'h0 : _GEN_935; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_937 = 10'h3a9 == index ? 32'h0 : _GEN_936; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_938 = 10'h3aa == index ? 32'h0 : _GEN_937; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_939 = 10'h3ab == index ? 32'h0 : _GEN_938; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_940 = 10'h3ac == index ? 32'h0 : _GEN_939; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_941 = 10'h3ad == index ? 32'h0 : _GEN_940; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_942 = 10'h3ae == index ? 32'h0 : _GEN_941; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_943 = 10'h3af == index ? 32'h0 : _GEN_942; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_944 = 10'h3b0 == index ? 32'h0 : _GEN_943; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_945 = 10'h3b1 == index ? 32'h0 : _GEN_944; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_946 = 10'h3b2 == index ? 32'h0 : _GEN_945; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_947 = 10'h3b3 == index ? 32'h0 : _GEN_946; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_948 = 10'h3b4 == index ? 32'h0 : _GEN_947; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_949 = 10'h3b5 == index ? 32'h0 : _GEN_948; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_950 = 10'h3b6 == index ? 32'h0 : _GEN_949; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_951 = 10'h3b7 == index ? 32'h0 : _GEN_950; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_952 = 10'h3b8 == index ? 32'h0 : _GEN_951; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_953 = 10'h3b9 == index ? 32'h0 : _GEN_952; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_954 = 10'h3ba == index ? 32'h0 : _GEN_953; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_955 = 10'h3bb == index ? 32'h0 : _GEN_954; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_956 = 10'h3bc == index ? 32'h0 : _GEN_955; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_957 = 10'h3bd == index ? 32'h0 : _GEN_956; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_958 = 10'h3be == index ? 32'h0 : _GEN_957; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_959 = 10'h3bf == index ? 32'h0 : _GEN_958; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_960 = 10'h3c0 == index ? 32'h0 : _GEN_959; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_961 = 10'h3c1 == index ? 32'h0 : _GEN_960; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_962 = 10'h3c2 == index ? 32'h0 : _GEN_961; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_963 = 10'h3c3 == index ? 32'h0 : _GEN_962; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_964 = 10'h3c4 == index ? 32'h0 : _GEN_963; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_965 = 10'h3c5 == index ? 32'h0 : _GEN_964; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_966 = 10'h3c6 == index ? 32'h0 : _GEN_965; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_967 = 10'h3c7 == index ? 32'h0 : _GEN_966; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_968 = 10'h3c8 == index ? 32'h0 : _GEN_967; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_969 = 10'h3c9 == index ? 32'h0 : _GEN_968; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_970 = 10'h3ca == index ? 32'h0 : _GEN_969; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_971 = 10'h3cb == index ? 32'h0 : _GEN_970; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_972 = 10'h3cc == index ? 32'h0 : _GEN_971; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_973 = 10'h3cd == index ? 32'h0 : _GEN_972; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_974 = 10'h3ce == index ? 32'h0 : _GEN_973; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_975 = 10'h3cf == index ? 32'h0 : _GEN_974; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_976 = 10'h3d0 == index ? 32'h0 : _GEN_975; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_977 = 10'h3d1 == index ? 32'h0 : _GEN_976; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_978 = 10'h3d2 == index ? 32'h0 : _GEN_977; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_979 = 10'h3d3 == index ? 32'h0 : _GEN_978; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_980 = 10'h3d4 == index ? 32'h0 : _GEN_979; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_981 = 10'h3d5 == index ? 32'h0 : _GEN_980; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_982 = 10'h3d6 == index ? 32'h0 : _GEN_981; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_983 = 10'h3d7 == index ? 32'h0 : _GEN_982; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_984 = 10'h3d8 == index ? 32'h0 : _GEN_983; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_985 = 10'h3d9 == index ? 32'h0 : _GEN_984; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_986 = 10'h3da == index ? 32'h0 : _GEN_985; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_987 = 10'h3db == index ? 32'h0 : _GEN_986; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_988 = 10'h3dc == index ? 32'h0 : _GEN_987; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_989 = 10'h3dd == index ? 32'h0 : _GEN_988; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_990 = 10'h3de == index ? 32'h0 : _GEN_989; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_991 = 10'h3df == index ? 32'h0 : _GEN_990; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_992 = 10'h3e0 == index ? 32'h0 : _GEN_991; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_993 = 10'h3e1 == index ? 32'h0 : _GEN_992; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_994 = 10'h3e2 == index ? 32'h0 : _GEN_993; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_995 = 10'h3e3 == index ? 32'h0 : _GEN_994; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_996 = 10'h3e4 == index ? 32'h0 : _GEN_995; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_997 = 10'h3e5 == index ? 32'h0 : _GEN_996; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_998 = 10'h3e6 == index ? 32'h0 : _GEN_997; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_999 = 10'h3e7 == index ? 32'h0 : _GEN_998; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1000 = 10'h3e8 == index ? 32'h0 : _GEN_999; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1001 = 10'h3e9 == index ? 32'h0 : _GEN_1000; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1002 = 10'h3ea == index ? 32'h0 : _GEN_1001; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1003 = 10'h3eb == index ? 32'h0 : _GEN_1002; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1004 = 10'h3ec == index ? 32'h0 : _GEN_1003; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1005 = 10'h3ed == index ? 32'h0 : _GEN_1004; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1006 = 10'h3ee == index ? 32'h0 : _GEN_1005; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1007 = 10'h3ef == index ? 32'h0 : _GEN_1006; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1008 = 10'h3f0 == index ? 32'h0 : _GEN_1007; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1009 = 10'h3f1 == index ? 32'h0 : _GEN_1008; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1010 = 10'h3f2 == index ? 32'h0 : _GEN_1009; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1011 = 10'h3f3 == index ? 32'h0 : _GEN_1010; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1012 = 10'h3f4 == index ? 32'h0 : _GEN_1011; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1013 = 10'h3f5 == index ? 32'h0 : _GEN_1012; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1014 = 10'h3f6 == index ? 32'h0 : _GEN_1013; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1015 = 10'h3f7 == index ? 32'h0 : _GEN_1014; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1016 = 10'h3f8 == index ? 32'h0 : _GEN_1015; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1017 = 10'h3f9 == index ? 32'h0 : _GEN_1016; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1018 = 10'h3fa == index ? 32'h0 : _GEN_1017; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1019 = 10'h3fb == index ? 32'h0 : _GEN_1018; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1020 = 10'h3fc == index ? 32'h0 : _GEN_1019; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1021 = 10'h3fd == index ? 32'h0 : _GEN_1020; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1022 = 10'h3fe == index ? 32'h0 : _GEN_1021; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign _GEN_1023 = 10'h3ff == index ? 32'h0 : _GEN_1022; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultRV32Config.fir@196968.4]
  assign auto_in_a_ready = auto_in_d_ready; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultRV32Config.fir@195936.4]
  assign auto_in_d_valid = auto_in_a_valid; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultRV32Config.fir@195936.4]
  assign auto_in_d_bits_size = auto_in_a_bits_size; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultRV32Config.fir@195936.4]
  assign auto_in_d_bits_source = auto_in_a_bits_source; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultRV32Config.fir@195936.4]
  assign auto_in_d_bits_data = _T ? 32'h0 : _GEN_1023; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultRV32Config.fir@195936.4]
  assign TLMonitor_clock = clock; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195914.4]
  assign TLMonitor_reset = reset; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@195915.4]
  assign TLMonitor_io_in_a_ready = auto_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195935.4]
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195934.4]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195933.4]
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195932.4]
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195931.4]
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195930.4]
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195929.4]
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195928.4]
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195926.4]
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195925.4]
  assign TLMonitor_io_in_d_valid = auto_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195924.4]
  assign TLMonitor_io_in_d_bits_size = auto_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195921.4]
  assign TLMonitor_io_in_d_bits_source = auto_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultRV32Config.fir@195920.4]
endmodule
