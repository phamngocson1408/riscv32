`include "include_module.v"
`ifdef __TLB
module TLB( 
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [31:0] io_req_bits_vaddr,
  input         io_req_bits_passthrough,
  input  [1:0]  io_req_bits_size, 
  input  [4:0]  io_req_bits_cmd,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_ld,
  output        io_resp_pf_st,
  output        io_resp_ae_ld,
  output        io_resp_ae_st,
  output        io_resp_ma_ld,
  output        io_resp_ma_st,
  output        io_resp_cacheable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [31:0] io_sfence_bits_addr,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [19:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn, 
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input         io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input         io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr, 
  input  [31:0] io_ptw_pmp_0_mask, 
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr, 
  input  [31:0] io_ptw_pmp_1_mask, 
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr, 
  input  [31:0] io_ptw_pmp_2_mask, 
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr, 
  input  [31:0] io_ptw_pmp_3_mask, 
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr, 
  input  [31:0] io_ptw_pmp_4_mask, 
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr, 
  input  [31:0] io_ptw_pmp_5_mask, 
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr, 
  input  [31:0] io_ptw_pmp_6_mask, 
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr, 
  input  [31:0] io_ptw_pmp_7_mask 
);
  wire [19:0] _2_io_x_ppn;
  wire  _2_io_x_u;
  wire  _2_io_x_ae;
  wire  _2_io_x_sw;
  wire  _2_io_x_sx;
  wire  _2_io_x_sr;
  wire  _2_io_x_pw;
  wire  _2_io_x_px;
  wire  _2_io_x_pr;
  wire  _2_io_x_pal;
  wire  _2_io_x_paa;
  wire  _2_io_x_eff;
  wire  _2_io_x_c;
  wire [19:0] _2_io_y_ppn;
  wire  _2_io_y_u;
  wire  _2_io_y_ae;
  wire  _2_io_y_sw;
  wire  _2_io_y_sx;
  wire  _2_io_y_sr;
  wire  _2_io_y_pw;
  wire  _2_io_y_px;
  wire  _2_io_y_pr;
  wire  _2_io_y_pal;
  wire  _2_io_y_paa;
  wire  _2_io_y_eff;
  wire  _2_io_y_c;
  wire [1:0] pmp_io_prv;
  wire  pmp_io_pmp_0_cfg_l;
  wire [1:0] pmp_io_pmp_0_cfg_a; 
  wire  pmp_io_pmp_0_cfg_x;
  wire  pmp_io_pmp_0_cfg_w; 
  wire  pmp_io_pmp_0_cfg_r;
  wire [29:0] pmp_io_pmp_0_addr;
  wire [31:0] pmp_io_pmp_0_mask;
  wire  pmp_io_pmp_1_cfg_l;
  wire [1:0] pmp_io_pmp_1_cfg_a;
  wire  pmp_io_pmp_1_cfg_x; 
  wire  pmp_io_pmp_1_cfg_w;
  wire  pmp_io_pmp_1_cfg_r;
  wire [29:0] pmp_io_pmp_1_addr;
  wire [31:0] pmp_io_pmp_1_mask;
  wire  pmp_io_pmp_2_cfg_l;
  wire [1:0] pmp_io_pmp_2_cfg_a;
  wire  pmp_io_pmp_2_cfg_x;
  wire  pmp_io_pmp_2_cfg_w;
  wire  pmp_io_pmp_2_cfg_r;
  wire [29:0] pmp_io_pmp_2_addr;
  wire [31:0] pmp_io_pmp_2_mask;
  wire  pmp_io_pmp_3_cfg_l;
  wire [1:0] pmp_io_pmp_3_cfg_a;
  wire  pmp_io_pmp_3_cfg_x;
  wire  pmp_io_pmp_3_cfg_w;
  wire  pmp_io_pmp_3_cfg_r;
  wire [29:0] pmp_io_pmp_3_addr;
  wire [31:0] pmp_io_pmp_3_mask;
  wire  pmp_io_pmp_4_cfg_l;
  wire [1:0] pmp_io_pmp_4_cfg_a;
  wire  pmp_io_pmp_4_cfg_x;
  wire  pmp_io_pmp_4_cfg_w;
  wire  pmp_io_pmp_4_cfg_r; 
  wire [29:0] pmp_io_pmp_4_addr;
  wire [31:0] pmp_io_pmp_4_mask;
  wire  pmp_io_pmp_5_cfg_l;
  wire [1:0] pmp_io_pmp_5_cfg_a;
  wire  pmp_io_pmp_5_cfg_x;
  wire  pmp_io_pmp_5_cfg_w;
  wire  pmp_io_pmp_5_cfg_r;
  wire [29:0] pmp_io_pmp_5_addr;
  wire [31:0] pmp_io_pmp_5_mask;
  wire  pmp_io_pmp_6_cfg_l;
  wire [1:0] pmp_io_pmp_6_cfg_a;
  wire  pmp_io_pmp_6_cfg_x; 
  wire  pmp_io_pmp_6_cfg_w; 
  wire  pmp_io_pmp_6_cfg_r;
  wire [29:0] pmp_io_pmp_6_addr;
  wire [31:0] pmp_io_pmp_6_mask;
  wire  pmp_io_pmp_7_cfg_l; 
  wire [1:0] pmp_io_pmp_7_cfg_a;
  wire  pmp_io_pmp_7_cfg_x;
  wire  pmp_io_pmp_7_cfg_w;
  wire  pmp_io_pmp_7_cfg_r;
  wire [29:0] pmp_io_pmp_7_addr; 
  wire [31:0] pmp_io_pmp_7_mask;
  wire [31:0] pmp_io_addr;
  wire  pmp_io_r;
  wire  pmp_io_w;
  wire  pmp_io_x; 
  wire [19:0] _2_1_io_x_ppn;
  wire  _2_1_io_x_u; 
  wire  _2_1_io_x_ae;
  wire  _2_1_io_x_sw;
  wire  _2_1_io_x_sx;
  wire  _2_1_io_x_sr;
  wire  _2_1_io_x_pw;
  wire  _2_1_io_x_px;
  wire  _2_1_io_x_pr;
  wire  _2_1_io_x_pal;
  wire  _2_1_io_x_paa; 
  wire  _2_1_io_x_eff;
  wire  _2_1_io_x_c;
  wire [19:0] _2_1_io_y_ppn;
  wire  _2_1_io_y_u;
  wire  _2_1_io_y_ae;
  wire  _2_1_io_y_sw;
  wire  _2_1_io_y_sx;
  wire  _2_1_io_y_sr;
  wire  _2_1_io_y_pw;
  wire  _2_1_io_y_px;
  wire  _2_1_io_y_pr;
  wire  _2_1_io_y_pal;
  wire  _2_1_io_y_paa;
  wire  _2_1_io_y_eff;
  wire  _2_1_io_y_c;
  wire [19:0] _2_2_io_x_ppn;
  wire  _2_2_io_x_u;
  wire  _2_2_io_x_ae;
  wire  _2_2_io_x_sw;
  wire  _2_2_io_x_sx;
  wire  _2_2_io_x_sr;
  wire  _2_2_io_x_pw;
  wire  _2_2_io_x_px;
  wire  _2_2_io_x_pr;
  wire  _2_2_io_x_pal;
  wire  _2_2_io_x_paa;
  wire  _2_2_io_x_eff;
  wire  _2_2_io_x_c;
  wire [19:0] _2_2_io_y_ppn;
  wire  _2_2_io_y_u;
  wire  _2_2_io_y_ae;
  wire  _2_2_io_y_sw;
  wire  _2_2_io_y_sx;
  wire  _2_2_io_y_sr;
  wire  _2_2_io_y_pw;
  wire  _2_2_io_y_px;
  wire  _2_2_io_y_pr;
  wire  _2_2_io_y_pal;
  wire  _2_2_io_y_paa;
  wire  _2_2_io_y_eff;
  wire  _2_2_io_y_c;
  wire [19:0] _2_3_io_x_ppn;
  wire  _2_3_io_x_u;
  wire  _2_3_io_x_ae;
  wire  _2_3_io_x_sw;
  wire  _2_3_io_x_sx;
  wire  _2_3_io_x_sr;
  wire  _2_3_io_x_pw;
  wire  _2_3_io_x_px;
  wire  _2_3_io_x_pr;
  wire  _2_3_io_x_pal;
  wire  _2_3_io_x_paa;
  wire  _2_3_io_x_eff;
  wire  _2_3_io_x_c;
  wire [19:0] _2_3_io_y_ppn;
  wire  _2_3_io_y_u;
  wire  _2_3_io_y_ae;
  wire  _2_3_io_y_sw;
  wire  _2_3_io_y_sx;
  wire  _2_3_io_y_sr;
  wire  _2_3_io_y_pw;
  wire  _2_3_io_y_px;
  wire  _2_3_io_y_pr;
  wire  _2_3_io_y_pal;
  wire  _2_3_io_y_paa;
  wire  _2_3_io_y_eff;
  wire  _2_3_io_y_c;
  wire [19:0] _2_4_io_x_ppn;
  wire  _2_4_io_x_u;
  wire  _2_4_io_x_ae;
  wire  _2_4_io_x_sw;
  wire  _2_4_io_x_sx;
  wire  _2_4_io_x_sr;
  wire  _2_4_io_x_pw;
  wire  _2_4_io_x_px;
  wire  _2_4_io_x_pr;
  wire  _2_4_io_x_pal;
  wire  _2_4_io_x_paa;
  wire  _2_4_io_x_eff;
  wire  _2_4_io_x_c;
  wire [19:0] _2_4_io_y_ppn;
  wire  _2_4_io_y_u;
  wire  _2_4_io_y_ae;
  wire  _2_4_io_y_sw;
  wire  _2_4_io_y_sx;
  wire  _2_4_io_y_sr;
  wire  _2_4_io_y_pw;
  wire  _2_4_io_y_px;
  wire  _2_4_io_y_pr;
  wire  _2_4_io_y_pal;
  wire  _2_4_io_y_paa;
  wire  _2_4_io_y_eff;
  wire  _2_4_io_y_c;
  wire [19:0] _2_5_io_x_ppn;
  wire  _2_5_io_x_u;
  wire  _2_5_io_x_ae;
  wire  _2_5_io_x_sw;
  wire  _2_5_io_x_sx;
  wire  _2_5_io_x_sr;
  wire  _2_5_io_x_pw;
  wire  _2_5_io_x_px;
  wire  _2_5_io_x_pr;
  wire  _2_5_io_x_pal;
  wire  _2_5_io_x_paa;
  wire  _2_5_io_x_eff;
  wire  _2_5_io_x_c;
  wire [19:0] _2_5_io_y_ppn;
  wire  _2_5_io_y_u;
  wire  _2_5_io_y_ae;
  wire  _2_5_io_y_sw;
  wire  _2_5_io_y_sx;
  wire  _2_5_io_y_sr;
  wire  _2_5_io_y_pw;
  wire  _2_5_io_y_px;
  wire  _2_5_io_y_pr;
  wire  _2_5_io_y_pal;
  wire  _2_5_io_y_paa;
  wire  _2_5_io_y_eff;
  wire  _2_5_io_y_c;
  wire [19:0] _2_6_io_x_ppn;
  wire  _2_6_io_x_u;
  wire  _2_6_io_x_ae;
  wire  _2_6_io_x_sw;
  wire  _2_6_io_x_sx;
  wire  _2_6_io_x_sr;
  wire  _2_6_io_x_pw;
  wire  _2_6_io_x_px;
  wire  _2_6_io_x_pr;
  wire  _2_6_io_x_pal;
  wire  _2_6_io_x_paa;
  wire  _2_6_io_x_eff;
  wire  _2_6_io_x_c;
  wire [19:0] _2_6_io_y_ppn;
  wire  _2_6_io_y_u;
  wire  _2_6_io_y_ae;
  wire  _2_6_io_y_sw;
  wire  _2_6_io_y_sx;
  wire  _2_6_io_y_sr;
  wire  _2_6_io_y_pw;
  wire  _2_6_io_y_px;
  wire  _2_6_io_y_pr;
  wire  _2_6_io_y_pal;
  wire  _2_6_io_y_paa;
  wire  _2_6_io_y_eff;
  wire  _2_6_io_y_c;
  wire [19:0] _2_7_io_x_ppn;
  wire  _2_7_io_x_u;
  wire  _2_7_io_x_ae;
  wire  _2_7_io_x_sw;
  wire  _2_7_io_x_sx;
  wire  _2_7_io_x_sr;
  wire  _2_7_io_x_pw;
  wire  _2_7_io_x_px;
  wire  _2_7_io_x_pr;
  wire  _2_7_io_x_pal;
  wire  _2_7_io_x_paa;
  wire  _2_7_io_x_eff;
  wire  _2_7_io_x_c;
  wire [19:0] _2_7_io_y_ppn;
  wire  _2_7_io_y_u;
  wire  _2_7_io_y_ae;
  wire  _2_7_io_y_sw;
  wire  _2_7_io_y_sx;
  wire  _2_7_io_y_sr;
  wire  _2_7_io_y_pw;
  wire  _2_7_io_y_px;
  wire  _2_7_io_y_pr;
  wire  _2_7_io_y_pal;
  wire  _2_7_io_y_paa;
  wire  _2_7_io_y_eff;
  wire  _2_7_io_y_c;
  wire [19:0] _2_8_io_x_ppn;
  wire  _2_8_io_x_u;
  wire  _2_8_io_x_ae;
  wire  _2_8_io_x_sw;
  wire  _2_8_io_x_sx;
  wire  _2_8_io_x_sr;
  wire  _2_8_io_x_pw;
  wire  _2_8_io_x_px;
  wire  _2_8_io_x_pr;
  wire  _2_8_io_x_pal;
  wire  _2_8_io_x_paa;
  wire  _2_8_io_x_eff;
  wire  _2_8_io_x_c;
  wire [19:0] _2_8_io_y_ppn;
  wire  _2_8_io_y_u;
  wire  _2_8_io_y_ae;
  wire  _2_8_io_y_sw;
  wire  _2_8_io_y_sx;
  wire  _2_8_io_y_sr;
  wire  _2_8_io_y_pw;
  wire  _2_8_io_y_px;
  wire  _2_8_io_y_pr;
  wire  _2_8_io_y_pal;
  wire  _2_8_io_y_paa;
  wire  _2_8_io_y_eff;
  wire  _2_8_io_y_c;
  wire [19:0] _2_9_io_x_ppn;
  wire  _2_9_io_x_u;
  wire  _2_9_io_x_ae;
  wire  _2_9_io_x_sw;
  wire  _2_9_io_x_sx;
  wire  _2_9_io_x_sr;
  wire  _2_9_io_x_pw;
  wire  _2_9_io_x_px;
  wire  _2_9_io_x_pr;
  wire  _2_9_io_x_pal;
  wire  _2_9_io_x_paa; 
  wire  _2_9_io_x_eff;
  wire  _2_9_io_x_c;
  wire [19:0] _2_9_io_y_ppn;
  wire  _2_9_io_y_u;
  wire  _2_9_io_y_ae;
  wire  _2_9_io_y_sw;
  wire  _2_9_io_y_sx;
  wire  _2_9_io_y_sr;
  wire  _2_9_io_y_pw;
  wire  _2_9_io_y_px;
  wire  _2_9_io_y_pr;
  wire  _2_9_io_y_pal;
  wire  _2_9_io_y_paa;
  wire  _2_9_io_y_eff;
  wire  _2_9_io_y_c;
  wire [19:0] _2_10_io_x_ppn;
  wire  _2_10_io_x_u;
  wire  _2_10_io_x_ae;
  wire  _2_10_io_x_sw;
  wire  _2_10_io_x_sx;
  wire  _2_10_io_x_sr;
  wire  _2_10_io_x_pw;
  wire  _2_10_io_x_px;
  wire  _2_10_io_x_pr;
  wire  _2_10_io_x_pal;
  wire  _2_10_io_x_paa;
  wire  _2_10_io_x_eff;
  wire  _2_10_io_x_c; 
  wire [19:0] _2_10_io_y_ppn;
  wire  _2_10_io_y_u;
  wire  _2_10_io_y_ae;
  wire  _2_10_io_y_sw;
  wire  _2_10_io_y_sx;
  wire  _2_10_io_y_sr;
  wire  _2_10_io_y_pw;
  wire  _2_10_io_y_px;
  wire  _2_10_io_y_pr;
  wire  _2_10_io_y_pal;
  wire  _2_10_io_y_paa;
  wire  _2_10_io_y_eff;
  wire  _2_10_io_y_c;
  wire [19:0] _2_11_io_x_ppn;
  wire  _2_11_io_x_u;
  wire  _2_11_io_x_ae;
  wire  _2_11_io_x_sw;
  wire  _2_11_io_x_sx;
  wire  _2_11_io_x_sr;
  wire  _2_11_io_x_pw;
  wire  _2_11_io_x_px;
  wire  _2_11_io_x_pr;
  wire  _2_11_io_x_pal;
  wire  _2_11_io_x_paa;
  wire  _2_11_io_x_eff;
  wire  _2_11_io_x_c; 
  wire [19:0] _2_11_io_y_ppn;
  wire  _2_11_io_y_u;
  wire  _2_11_io_y_ae;
  wire  _2_11_io_y_sw;
  wire  _2_11_io_y_sx;
  wire  _2_11_io_y_sr;
  wire  _2_11_io_y_pw;
  wire  _2_11_io_y_px;
  wire  _2_11_io_y_pr;
  wire  _2_11_io_y_pal; 
  wire  _2_11_io_y_paa; 
  wire  _2_11_io_y_eff;
  wire  _2_11_io_y_c;
  wire [19:0] _2_12_io_x_ppn;
  wire  _2_12_io_x_u; 
  wire  _2_12_io_x_ae; 
  wire  _2_12_io_x_sw; 
  wire  _2_12_io_x_sx; 
  wire  _2_12_io_x_sr; 
  wire  _2_12_io_x_pw; 
  wire  _2_12_io_x_px; 
  wire  _2_12_io_x_pr; 
  wire  _2_12_io_x_pal;
  wire  _2_12_io_x_paa;
  wire  _2_12_io_x_eff;
  wire  _2_12_io_x_c;
  wire [19:0] _2_12_io_y_ppn;
  wire  _2_12_io_y_u; 
  wire  _2_12_io_y_ae;
  wire  _2_12_io_y_sw;
  wire  _2_12_io_y_sx;
  wire  _2_12_io_y_sr;
  wire  _2_12_io_y_pw;
  wire  _2_12_io_y_px;
  wire  _2_12_io_y_pr;
  wire  _2_12_io_y_pal;
  wire  _2_12_io_y_paa;
  wire  _2_12_io_y_eff;
  wire  _2_12_io_y_c;
  wire [19:0] _2_13_io_x_ppn;
  wire  _2_13_io_x_u;
  wire  _2_13_io_x_ae;
  wire  _2_13_io_x_sw;
  wire  _2_13_io_x_sx;
  wire  _2_13_io_x_sr;
  wire  _2_13_io_x_pw;
  wire  _2_13_io_x_px;
  wire  _2_13_io_x_pr;
  wire  _2_13_io_x_pal;
  wire  _2_13_io_x_paa;
  wire  _2_13_io_x_eff;
  wire  _2_13_io_x_c;
  wire [19:0] _2_13_io_y_ppn;
  wire  _2_13_io_y_u;
  wire  _2_13_io_y_ae;
  wire  _2_13_io_y_sw;
  wire  _2_13_io_y_sx;
  wire  _2_13_io_y_sr;
  wire  _2_13_io_y_pw;
  wire  _2_13_io_y_px;
  wire  _2_13_io_y_pr;
  wire  _2_13_io_y_pal;
  wire  _2_13_io_y_paa;
  wire  _2_13_io_y_eff;
  wire  _2_13_io_y_c;
  wire [19:0] _2_14_io_x_ppn;
  wire  _2_14_io_x_u;
  wire  _2_14_io_x_ae;
  wire  _2_14_io_x_sw;
  wire  _2_14_io_x_sx;
  wire  _2_14_io_x_sr;
  wire  _2_14_io_x_pw;
  wire  _2_14_io_x_px;
  wire  _2_14_io_x_pr;
  wire  _2_14_io_x_pal;
  wire  _2_14_io_x_paa;
  wire  _2_14_io_x_eff;
  wire  _2_14_io_x_c;
  wire [19:0] _2_14_io_y_ppn;
  wire  _2_14_io_y_u;
  wire  _2_14_io_y_ae;
  wire  _2_14_io_y_sw;
  wire  _2_14_io_y_sx;
  wire  _2_14_io_y_sr;
  wire  _2_14_io_y_pw;
  wire  _2_14_io_y_px;
  wire  _2_14_io_y_pr;
  wire  _2_14_io_y_pal;
  wire  _2_14_io_y_paa;
  wire  _2_14_io_y_eff;
  wire  _2_14_io_y_c;
  wire [19:0] _2_15_io_x_ppn;
  wire  _2_15_io_x_u;
  wire  _2_15_io_x_ae;
  wire  _2_15_io_x_sw;
  wire  _2_15_io_x_sx;
  wire  _2_15_io_x_sr;
  wire  _2_15_io_x_pw;
  wire  _2_15_io_x_px;
  wire  _2_15_io_x_pr;
  wire  _2_15_io_x_pal;
  wire  _2_15_io_x_paa; 
  wire  _2_15_io_x_eff;
  wire  _2_15_io_x_c;
  wire [19:0] _2_15_io_y_ppn;
  wire  _2_15_io_y_u;
  wire  _2_15_io_y_ae;
  wire  _2_15_io_y_sw;
  wire  _2_15_io_y_sx;
  wire  _2_15_io_y_sr;
  wire  _2_15_io_y_pw;
  wire  _2_15_io_y_px;
  wire  _2_15_io_y_pr;
  wire  _2_15_io_y_pal;
  wire  _2_15_io_y_paa;
  wire  _2_15_io_y_eff;
  wire  _2_15_io_y_c;
  wire [19:0] _2_16_io_x_ppn;
  wire  _2_16_io_x_u;
  wire  _2_16_io_x_ae;
  wire  _2_16_io_x_sw;
  wire  _2_16_io_x_sx;
  wire  _2_16_io_x_sr;
  wire  _2_16_io_x_pw;
  wire  _2_16_io_x_px;
  wire  _2_16_io_x_pr;
  wire  _2_16_io_x_pal;
  wire  _2_16_io_x_paa;
  wire  _2_16_io_x_eff;
  wire  _2_16_io_x_c;
  wire [19:0] _2_16_io_y_ppn;
  wire  _2_16_io_y_u;
  wire  _2_16_io_y_ae;
  wire  _2_16_io_y_sw;
  wire  _2_16_io_y_sx;
  wire  _2_16_io_y_sr;
  wire  _2_16_io_y_pw;
  wire  _2_16_io_y_px;
  wire  _2_16_io_y_pr;
  wire  _2_16_io_y_pal;
  wire  _2_16_io_y_paa;
  wire  _2_16_io_y_eff; 
  wire  _2_16_io_y_c;
  wire [19:0] _2_17_io_x_ppn;
  wire  _2_17_io_x_u;
  wire  _2_17_io_x_ae;
  wire  _2_17_io_x_sw;
  wire  _2_17_io_x_sx;
  wire  _2_17_io_x_sr;
  wire  _2_17_io_x_pw;
  wire  _2_17_io_x_px;
  wire  _2_17_io_x_pr;
  wire  _2_17_io_x_pal;
  wire  _2_17_io_x_paa;
  wire  _2_17_io_x_eff;
  wire  _2_17_io_x_c;
  wire [19:0] _2_17_io_y_ppn;
  wire  _2_17_io_y_u;
  wire  _2_17_io_y_ae;
  wire  _2_17_io_y_sw;
  wire  _2_17_io_y_sx;
  wire  _2_17_io_y_sr;
  wire  _2_17_io_y_pw;
  wire  _2_17_io_y_px;
  wire  _2_17_io_y_pr;
  wire  _2_17_io_y_pal;
  wire  _2_17_io_y_paa;
  wire  _2_17_io_y_eff;
  wire  _2_17_io_y_c;
  wire [19:0] _2_18_io_x_ppn;
  wire  _2_18_io_x_u;
  wire  _2_18_io_x_ae;
  wire  _2_18_io_x_sw;
  wire  _2_18_io_x_sx;
  wire  _2_18_io_x_sr;
  wire  _2_18_io_x_pw;
  wire  _2_18_io_x_px;
  wire  _2_18_io_x_pr;
  wire  _2_18_io_x_pal;
  wire  _2_18_io_x_paa;
  wire  _2_18_io_x_eff;
  wire  _2_18_io_x_c;
  wire [19:0] _2_18_io_y_ppn;
  wire  _2_18_io_y_u;
  wire  _2_18_io_y_ae;
  wire  _2_18_io_y_sw;
  wire  _2_18_io_y_sx;
  wire  _2_18_io_y_sr;
  wire  _2_18_io_y_pw;
  wire  _2_18_io_y_px;
  wire  _2_18_io_y_pr;
  wire  _2_18_io_y_pal;
  wire  _2_18_io_y_paa;
  wire  _2_18_io_y_eff;
  wire  _2_18_io_y_c;
  wire [19:0] _2_19_io_x_ppn;
  wire  _2_19_io_x_u;
  wire  _2_19_io_x_ae;
  wire  _2_19_io_x_sw;
  wire  _2_19_io_x_sx;
  wire  _2_19_io_x_sr;
  wire  _2_19_io_x_pw;
  wire  _2_19_io_x_px;
  wire  _2_19_io_x_pr;
  wire  _2_19_io_x_pal;
  wire  _2_19_io_x_paa; 
  wire  _2_19_io_x_eff;
  wire  _2_19_io_x_c;
  wire [19:0] _2_19_io_y_ppn;
  wire  _2_19_io_y_u;
  wire  _2_19_io_y_ae;
  wire  _2_19_io_y_sw;
  wire  _2_19_io_y_sx;
  wire  _2_19_io_y_sr;
  wire  _2_19_io_y_pw;
  wire  _2_19_io_y_px;
  wire  _2_19_io_y_pr;
  wire  _2_19_io_y_pal;
  wire  _2_19_io_y_paa;
  wire  _2_19_io_y_eff;
  wire  _2_19_io_y_c;
  wire [19:0] _2_20_io_x_ppn;
  wire  _2_20_io_x_u;
  wire  _2_20_io_x_ae;
  wire  _2_20_io_x_sw;
  wire  _2_20_io_x_sx;
  wire  _2_20_io_x_sr;
  wire  _2_20_io_x_pw;
  wire  _2_20_io_x_px;
  wire  _2_20_io_x_pr;
  wire  _2_20_io_x_pal;
  wire  _2_20_io_x_paa;
  wire  _2_20_io_x_eff;
  wire  _2_20_io_x_c;
  wire [19:0] _2_20_io_y_ppn;
  wire  _2_20_io_y_u;
  wire  _2_20_io_y_ae;
  wire  _2_20_io_y_sw;
  wire  _2_20_io_y_sx;
  wire  _2_20_io_y_sr;
  wire  _2_20_io_y_pw;
  wire  _2_20_io_y_px;
  wire  _2_20_io_y_pr;
  wire  _2_20_io_y_pal;
  wire  _2_20_io_y_paa;
  wire  _2_20_io_y_eff;
  wire  _2_20_io_y_c;
  wire [19:0] _2_21_io_x_ppn;
  wire  _2_21_io_x_u;
  wire  _2_21_io_x_ae;
  wire  _2_21_io_x_sw;
  wire  _2_21_io_x_sx;
  wire  _2_21_io_x_sr;
  wire  _2_21_io_x_pw;
  wire  _2_21_io_x_px;
  wire  _2_21_io_x_pr;
  wire  _2_21_io_x_pal;
  wire  _2_21_io_x_paa;
  wire  _2_21_io_x_eff;
  wire  _2_21_io_x_c;
  wire [19:0] _2_21_io_y_ppn;
  wire  _2_21_io_y_u;
  wire  _2_21_io_y_ae;
  wire  _2_21_io_y_sw;
  wire  _2_21_io_y_sx;
  wire  _2_21_io_y_sr;
  wire  _2_21_io_y_pw;
  wire  _2_21_io_y_px;
  wire  _2_21_io_y_pr;
  wire  _2_21_io_y_pal;
  wire  _2_21_io_y_paa;
  wire  _2_21_io_y_eff;
  wire  _2_21_io_y_c;
  wire [19:0] _2_22_io_x_ppn;
  wire  _2_22_io_x_u;
  wire  _2_22_io_x_ae;
  wire  _2_22_io_x_sw;
  wire  _2_22_io_x_sx;
  wire  _2_22_io_x_sr;
  wire  _2_22_io_x_pw;
  wire  _2_22_io_x_px;
  wire  _2_22_io_x_pr;
  wire  _2_22_io_x_pal;
  wire  _2_22_io_x_paa;
  wire  _2_22_io_x_eff;
  wire  _2_22_io_x_c;
  wire [19:0] _2_22_io_y_ppn;
  wire  _2_22_io_y_u;
  wire  _2_22_io_y_ae;
  wire  _2_22_io_y_sw;
  wire  _2_22_io_y_sx;
  wire  _2_22_io_y_sr;
  wire  _2_22_io_y_pw;
  wire  _2_22_io_y_px;
  wire  _2_22_io_y_pr;
  wire  _2_22_io_y_pal;
  wire  _2_22_io_y_paa;
  wire  _2_22_io_y_eff;
  wire  _2_22_io_y_c;
  wire [19:0] _2_23_io_x_ppn; 
  wire  _2_23_io_x_u;
  wire  _2_23_io_x_ae;
  wire  _2_23_io_x_sw;
  wire  _2_23_io_x_sx;
  wire  _2_23_io_x_sr;
  wire  _2_23_io_x_pw;
  wire  _2_23_io_x_px;
  wire  _2_23_io_x_pr;
  wire  _2_23_io_x_pal;
  wire  _2_23_io_x_paa;
  wire  _2_23_io_x_eff;
  wire  _2_23_io_x_c;
  wire [19:0] _2_23_io_y_ppn;
  wire  _2_23_io_y_u;
  wire  _2_23_io_y_ae;
  wire  _2_23_io_y_sw;
  wire  _2_23_io_y_sx;
  wire  _2_23_io_y_sr;
  wire  _2_23_io_y_pw;
  wire  _2_23_io_y_px;
  wire  _2_23_io_y_pr;
  wire  _2_23_io_y_pal;
  wire  _2_23_io_y_paa;
  wire  _2_23_io_y_eff;
  wire  _2_23_io_y_c;
  wire [19:0] _2_24_io_x_ppn;
  wire  _2_24_io_x_u;
  wire  _2_24_io_x_ae;
  wire  _2_24_io_x_sw;
  wire  _2_24_io_x_sx;
  wire  _2_24_io_x_sr;
  wire  _2_24_io_x_pw;
  wire  _2_24_io_x_px;
  wire  _2_24_io_x_pr;
  wire  _2_24_io_x_pal;
  wire  _2_24_io_x_paa;
  wire  _2_24_io_x_eff;
  wire  _2_24_io_x_c;
  wire [19:0] _2_24_io_y_ppn;
  wire  _2_24_io_y_u;
  wire  _2_24_io_y_ae;
  wire  _2_24_io_y_sw;
  wire  _2_24_io_y_sx;
  wire  _2_24_io_y_sr;
  wire  _2_24_io_y_pw;
  wire  _2_24_io_y_px;
  wire  _2_24_io_y_pr;
  wire  _2_24_io_y_pal;
  wire  _2_24_io_y_paa;
  wire  _2_24_io_y_eff;
  wire  _2_24_io_y_c;
  wire [19:0] _2_25_io_x_ppn;
  wire  _2_25_io_x_u;
  wire  _2_25_io_x_ae;
  wire  _2_25_io_x_sw;
  wire  _2_25_io_x_sx;
  wire  _2_25_io_x_sr;
  wire  _2_25_io_x_pw;
  wire  _2_25_io_x_px;
  wire  _2_25_io_x_pr;
  wire  _2_25_io_x_pal;
  wire  _2_25_io_x_paa;
  wire  _2_25_io_x_eff;
  wire  _2_25_io_x_c;
  wire [19:0] _2_25_io_y_ppn;
  wire  _2_25_io_y_u;
  wire  _2_25_io_y_ae;
  wire  _2_25_io_y_sw;
  wire  _2_25_io_y_sx;
  wire  _2_25_io_y_sr;
  wire  _2_25_io_y_pw;
  wire  _2_25_io_y_px;
  wire  _2_25_io_y_pr;
  wire  _2_25_io_y_pal;
  wire  _2_25_io_y_paa;
  wire  _2_25_io_y_eff;
  wire  _2_25_io_y_c;
  wire [19:0] _2_26_io_x_ppn;
  wire  _2_26_io_x_u;
  wire  _2_26_io_x_ae;
  wire  _2_26_io_x_sw;
  wire  _2_26_io_x_sx;
  wire  _2_26_io_x_sr;
  wire  _2_26_io_x_pw;
  wire  _2_26_io_x_px;
  wire  _2_26_io_x_pr;
  wire  _2_26_io_x_pal;
  wire  _2_26_io_x_paa;
  wire  _2_26_io_x_eff;
  wire  _2_26_io_x_c;
  wire [19:0] _2_26_io_y_ppn;
  wire  _2_26_io_y_u;
  wire  _2_26_io_y_ae;
  wire  _2_26_io_y_sw;
  wire  _2_26_io_y_sx;
  wire  _2_26_io_y_sr;
  wire  _2_26_io_y_pw;
  wire  _2_26_io_y_px;
  wire  _2_26_io_y_pr;
  wire  _2_26_io_y_pal;
  wire  _2_26_io_y_paa;
  wire  _2_26_io_y_eff;
  wire  _2_26_io_y_c;
  wire [19:0] _2_27_io_x_ppn;
  wire  _2_27_io_x_u;
  wire  _2_27_io_x_ae;
  wire  _2_27_io_x_sw;
  wire  _2_27_io_x_sx;
  wire  _2_27_io_x_sr;
  wire  _2_27_io_x_pw;
  wire  _2_27_io_x_px;
  wire  _2_27_io_x_pr;
  wire  _2_27_io_x_pal;
  wire  _2_27_io_x_paa;
  wire  _2_27_io_x_eff;
  wire  _2_27_io_x_c;
  wire [19:0] _2_27_io_y_ppn;
  wire  _2_27_io_y_u;
  wire  _2_27_io_y_ae;
  wire  _2_27_io_y_sw;
  wire  _2_27_io_y_sx;
  wire  _2_27_io_y_sr;
  wire  _2_27_io_y_pw;
  wire  _2_27_io_y_px;
  wire  _2_27_io_y_pr;
  wire  _2_27_io_y_pal;
  wire  _2_27_io_y_paa;
  wire  _2_27_io_y_eff;
  wire  _2_27_io_y_c;
  wire [19:0] _2_28_io_x_ppn;
  wire  _2_28_io_x_u;
  wire  _2_28_io_x_ae;
  wire  _2_28_io_x_sw;
  wire  _2_28_io_x_sx;
  wire  _2_28_io_x_sr;
  wire  _2_28_io_x_pw;
  wire  _2_28_io_x_px;
  wire  _2_28_io_x_pr;
  wire  _2_28_io_x_pal;
  wire  _2_28_io_x_paa;
  wire  _2_28_io_x_eff;
  wire  _2_28_io_x_c;
  wire [19:0] _2_28_io_y_ppn;
  wire  _2_28_io_y_u;
  wire  _2_28_io_y_ae;
  wire  _2_28_io_y_sw;
  wire  _2_28_io_y_sx;
  wire  _2_28_io_y_sr;
  wire  _2_28_io_y_pw;
  wire  _2_28_io_y_px;
  wire  _2_28_io_y_pr;
  wire  _2_28_io_y_pal;
  wire  _2_28_io_y_paa;
  wire  _2_28_io_y_eff; 
  wire  _2_28_io_y_c;
  wire [19:0] _2_29_io_x_ppn;
  wire  _2_29_io_x_u;
  wire  _2_29_io_x_ae;
  wire  _2_29_io_x_sw;
  wire  _2_29_io_x_sx;
  wire  _2_29_io_x_sr;
  wire  _2_29_io_x_pw;
  wire  _2_29_io_x_px;
  wire  _2_29_io_x_pr;
  wire  _2_29_io_x_pal;
  wire  _2_29_io_x_paa;
  wire  _2_29_io_x_eff;
  wire  _2_29_io_x_c;
  wire [19:0] _2_29_io_y_ppn;
  wire  _2_29_io_y_u;
  wire  _2_29_io_y_ae;
  wire  _2_29_io_y_sw;
  wire  _2_29_io_y_sx;
  wire  _2_29_io_y_sr;
  wire  _2_29_io_y_pw;
  wire  _2_29_io_y_px;
  wire  _2_29_io_y_pr;
  wire  _2_29_io_y_pal;
  wire  _2_29_io_y_paa;
  wire  _2_29_io_y_eff;
  wire  _2_29_io_y_c;
  wire [19:0] _2_30_io_x_ppn;
  wire  _2_30_io_x_u;
  wire  _2_30_io_x_ae;
  wire  _2_30_io_x_sw;
  wire  _2_30_io_x_sx;
  wire  _2_30_io_x_sr;
  wire  _2_30_io_x_pw;
  wire  _2_30_io_x_px;
  wire  _2_30_io_x_pr;
  wire  _2_30_io_x_pal;
  wire  _2_30_io_x_paa;
  wire  _2_30_io_x_eff;
  wire  _2_30_io_x_c;
  wire [19:0] _2_30_io_y_ppn;
  wire  _2_30_io_y_u;
  wire  _2_30_io_y_ae;
  wire  _2_30_io_y_sw;
  wire  _2_30_io_y_sx;
  wire  _2_30_io_y_sr;
  wire  _2_30_io_y_pw;
  wire  _2_30_io_y_px;
  wire  _2_30_io_y_pr;
  wire  _2_30_io_y_pal;
  wire  _2_30_io_y_paa; 
  wire  _2_30_io_y_eff;
  wire  _2_30_io_y_c; 
  wire [19:0] _2_31_io_x_ppn;
  wire  _2_31_io_x_u;
  wire  _2_31_io_x_ae;
  wire  _2_31_io_x_sw;
  wire  _2_31_io_x_sx;
  wire  _2_31_io_x_sr;
  wire  _2_31_io_x_pw;
  wire  _2_31_io_x_px;
  wire  _2_31_io_x_pr;
  wire  _2_31_io_x_pal;
  wire  _2_31_io_x_paa; 
  wire  _2_31_io_x_eff;
  wire  _2_31_io_x_c;
  wire [19:0] _2_31_io_y_ppn;
  wire  _2_31_io_y_u;
  wire  _2_31_io_y_ae;
  wire  _2_31_io_y_sw;
  wire  _2_31_io_y_sx;
  wire  _2_31_io_y_sr;
  wire  _2_31_io_y_pw;
  wire  _2_31_io_y_px;
  wire  _2_31_io_y_pr;
  wire  _2_31_io_y_pal;
  wire  _2_31_io_y_paa; 
  wire  _2_31_io_y_eff;
  wire  _2_31_io_y_c;
  wire [19:0] _2_32_io_x_ppn;
  wire  _2_32_io_x_u;
  wire  _2_32_io_x_ae;
  wire  _2_32_io_x_sw;
  wire  _2_32_io_x_sx;
  wire  _2_32_io_x_sr;
  wire  _2_32_io_x_pw;
  wire  _2_32_io_x_px;
  wire  _2_32_io_x_pr;
  wire  _2_32_io_x_pal;
  wire  _2_32_io_x_paa;
  wire  _2_32_io_x_eff;
  wire  _2_32_io_x_c;
  wire [19:0] _2_32_io_y_ppn;
  wire  _2_32_io_y_u;
  wire  _2_32_io_y_ae;
  wire  _2_32_io_y_sw;
  wire  _2_32_io_y_sx;
  wire  _2_32_io_y_sr;
  wire  _2_32_io_y_pw;
  wire  _2_32_io_y_px;
  wire  _2_32_io_y_pr;
  wire  _2_32_io_y_pal;
  wire  _2_32_io_y_paa;
  wire  _2_32_io_y_eff;
  wire  _2_32_io_y_c;
  wire [19:0] _2_33_io_x_ppn;
  wire  _2_33_io_x_u;
  wire  _2_33_io_x_ae;
  wire  _2_33_io_x_sw;
  wire  _2_33_io_x_sx;
  wire  _2_33_io_x_sr;
  wire  _2_33_io_x_pw;
  wire  _2_33_io_x_px;
  wire  _2_33_io_x_pr;
  wire  _2_33_io_x_pal;
  wire  _2_33_io_x_paa;
  wire  _2_33_io_x_eff;
  wire  _2_33_io_x_c;
  wire [19:0] _2_33_io_y_ppn;
  wire  _2_33_io_y_u; 
  wire  _2_33_io_y_ae;
  wire  _2_33_io_y_sw;
  wire  _2_33_io_y_sx;
  wire  _2_33_io_y_sr;
  wire  _2_33_io_y_pw;
  wire  _2_33_io_y_px;
  wire  _2_33_io_y_pr;
  wire  _2_33_io_y_pal;
  wire  _2_33_io_y_paa;
  wire  _2_33_io_y_eff;
  wire  _2_33_io_y_c;
  wire [19:0] _2_34_io_x_ppn;
  wire  _2_34_io_x_u;
  wire  _2_34_io_x_ae;
  wire  _2_34_io_x_sw;
  wire  _2_34_io_x_sx;
  wire  _2_34_io_x_sr;
  wire  _2_34_io_x_pw;
  wire  _2_34_io_x_px;
  wire  _2_34_io_x_pr;
  wire  _2_34_io_x_pal;
  wire  _2_34_io_x_paa;
  wire  _2_34_io_x_eff;
  wire  _2_34_io_x_c;
  wire [19:0] _2_34_io_y_ppn;
  wire  _2_34_io_y_u;
  wire  _2_34_io_y_ae;
  wire  _2_34_io_y_sw;
  wire  _2_34_io_y_sx;
  wire  _2_34_io_y_sr;
  wire  _2_34_io_y_pw;
  wire  _2_34_io_y_px;
  wire  _2_34_io_y_pr;
  wire  _2_34_io_y_pal;
  wire  _2_34_io_y_paa;
  wire  _2_34_io_y_eff;
  wire  _2_34_io_y_c;
  wire [19:0] _2_35_io_x_ppn;
  wire  _2_35_io_x_u;
  wire  _2_35_io_x_ae;
  wire  _2_35_io_x_sw;
  wire  _2_35_io_x_sx;
  wire  _2_35_io_x_sr;
  wire  _2_35_io_x_pw;
  wire  _2_35_io_x_px;
  wire  _2_35_io_x_pr;
  wire  _2_35_io_x_pal;
  wire  _2_35_io_x_paa;
  wire  _2_35_io_x_eff;
  wire  _2_35_io_x_c;
  wire [19:0] _2_35_io_y_ppn;
  wire  _2_35_io_y_u;
  wire  _2_35_io_y_ae;
  wire  _2_35_io_y_sw;
  wire  _2_35_io_y_sx;
  wire  _2_35_io_y_sr;
  wire  _2_35_io_y_pw;
  wire  _2_35_io_y_px;
  wire  _2_35_io_y_pr;
  wire  _2_35_io_y_pal;
  wire  _2_35_io_y_paa;
  wire  _2_35_io_y_eff;
  wire  _2_35_io_y_c;
  wire [19:0] _2_36_io_x_ppn;
  wire  _2_36_io_x_u;
  wire  _2_36_io_x_ae;
  wire  _2_36_io_x_sw;
  wire  _2_36_io_x_sx;
  wire  _2_36_io_x_sr;
  wire  _2_36_io_x_pw;
  wire  _2_36_io_x_px;
  wire  _2_36_io_x_pr;
  wire  _2_36_io_x_pal;
  wire  _2_36_io_x_paa;
  wire  _2_36_io_x_eff;
  wire  _2_36_io_x_c;
  wire [19:0] _2_36_io_y_ppn;
  wire  _2_36_io_y_u;
  wire  _2_36_io_y_ae;
  wire  _2_36_io_y_sw;
  wire  _2_36_io_y_sx;
  wire  _2_36_io_y_sr;
  wire  _2_36_io_y_pw;
  wire  _2_36_io_y_px;
  wire  _2_36_io_y_pr;
  wire  _2_36_io_y_pal;
  wire  _2_36_io_y_paa;
  wire  _2_36_io_y_eff;
  wire  _2_36_io_y_c;
  wire [19:0] _2_37_io_x_ppn;
  wire  _2_37_io_x_u;
  wire  _2_37_io_x_ae;
  wire  _2_37_io_x_sw;
  wire  _2_37_io_x_sx;
  wire  _2_37_io_x_sr;
  wire  _2_37_io_x_pw;
  wire  _2_37_io_x_px;
  wire  _2_37_io_x_pr;
  wire  _2_37_io_x_pal;
  wire  _2_37_io_x_paa;
  wire  _2_37_io_x_eff;
  wire  _2_37_io_x_c;
  wire [19:0] _2_37_io_y_ppn;
  wire  _2_37_io_y_u;
  wire  _2_37_io_y_ae;
  wire  _2_37_io_y_sw;
  wire  _2_37_io_y_sx;
  wire  _2_37_io_y_sr;
  wire  _2_37_io_y_pw;
  wire  _2_37_io_y_px;
  wire  _2_37_io_y_pr;
  wire  _2_37_io_y_pal;
  wire  _2_37_io_y_paa;
  wire  _2_37_io_y_eff;
  wire  _2_37_io_y_c;
  wire [19:0] _2_38_io_x_ppn;
  wire  _2_38_io_x_u;
  wire  _2_38_io_x_ae;
  wire  _2_38_io_x_sw;
  wire  _2_38_io_x_sx;
  wire  _2_38_io_x_sr;
  wire  _2_38_io_x_pw;
  wire  _2_38_io_x_px;
  wire  _2_38_io_x_pr;
  wire  _2_38_io_x_pal;
  wire  _2_38_io_x_paa;
  wire  _2_38_io_x_eff;
  wire  _2_38_io_x_c;
  wire [19:0] _2_38_io_y_ppn;
  wire  _2_38_io_y_u;
  wire  _2_38_io_y_ae;
  wire  _2_38_io_y_sw;
  wire  _2_38_io_y_sx;
  wire  _2_38_io_y_sr;
  wire  _2_38_io_y_pw;
  wire  _2_38_io_y_px;
  wire  _2_38_io_y_pr;
  wire  _2_38_io_y_pal;
  wire  _2_38_io_y_paa;
  wire  _2_38_io_y_eff;
  wire  _2_38_io_y_c;
  reg [19:0] sectored_entries_0_tag;
  reg [31:0] _RAND_0;
  reg [33:0] sectored_entries_0_data_0;
  reg [63:0] _RAND_1;
  reg [33:0] sectored_entries_0_data_1; 
  reg [63:0] _RAND_2;
  reg [33:0] sectored_entries_0_data_2; 
  reg [63:0] _RAND_3;
  reg [33:0] sectored_entries_0_data_3;
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_valid_0;
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_valid_1;
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_valid_2;
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_valid_3;
  reg [31:0] _RAND_8;
  reg [19:0] sectored_entries_1_tag; 
  reg [31:0] _RAND_9;
  reg [33:0] sectored_entries_1_data_0;
  reg [63:0] _RAND_10;
  reg [33:0] sectored_entries_1_data_1;
  reg [63:0] _RAND_11;
  reg [33:0] sectored_entries_1_data_2; 
  reg [63:0] _RAND_12;
  reg [33:0] sectored_entries_1_data_3; 
  reg [63:0] _RAND_13;
  reg  sectored_entries_1_valid_0;
  reg [31:0] _RAND_14;
  reg  sectored_entries_1_valid_1; 
  reg [31:0] _RAND_15;
  reg  sectored_entries_1_valid_2;
  reg [31:0] _RAND_16;
  reg  sectored_entries_1_valid_3;
  reg [31:0] _RAND_17;
  reg [19:0] sectored_entries_2_tag;
  reg [31:0] _RAND_18;
  reg [33:0] sectored_entries_2_data_0;
  reg [63:0] _RAND_19;
  reg [33:0] sectored_entries_2_data_1;
  reg [63:0] _RAND_20;
  reg [33:0] sectored_entries_2_data_2;
  reg [63:0] _RAND_21;
  reg [33:0] sectored_entries_2_data_3;
  reg [63:0] _RAND_22;
  reg  sectored_entries_2_valid_0;
  reg [31:0] _RAND_23;
  reg  sectored_entries_2_valid_1;
  reg [31:0] _RAND_24;
  reg  sectored_entries_2_valid_2;
  reg [31:0] _RAND_25;
  reg  sectored_entries_2_valid_3;
  reg [31:0] _RAND_26;
  reg [19:0] sectored_entries_3_tag;
  reg [31:0] _RAND_27;
  reg [33:0] sectored_entries_3_data_0;
  reg [63:0] _RAND_28;
  reg [33:0] sectored_entries_3_data_1;
  reg [63:0] _RAND_29;
  reg [33:0] sectored_entries_3_data_2;
  reg [63:0] _RAND_30;
  reg [33:0] sectored_entries_3_data_3;
  reg [63:0] _RAND_31;
  reg  sectored_entries_3_valid_0; 
  reg [31:0] _RAND_32;
  reg  sectored_entries_3_valid_1; 
  reg [31:0] _RAND_33;
  reg  sectored_entries_3_valid_2; 
  reg [31:0] _RAND_34;
  reg  sectored_entries_3_valid_3; 
  reg [31:0] _RAND_35;
  reg [19:0] sectored_entries_4_tag;
  reg [31:0] _RAND_36;
  reg [33:0] sectored_entries_4_data_0; 
  reg [63:0] _RAND_37;
  reg [33:0] sectored_entries_4_data_1;
  reg [63:0] _RAND_38;
  reg [33:0] sectored_entries_4_data_2;
  reg [63:0] _RAND_39;
  reg [33:0] sectored_entries_4_data_3;
  reg [63:0] _RAND_40;
  reg  sectored_entries_4_valid_0;
  reg [31:0] _RAND_41;
  reg  sectored_entries_4_valid_1;
  reg [31:0] _RAND_42;
  reg  sectored_entries_4_valid_2;
  reg [31:0] _RAND_43;
  reg  sectored_entries_4_valid_3;
  reg [31:0] _RAND_44;
  reg [19:0] sectored_entries_5_tag;
  reg [31:0] _RAND_45;
  reg [33:0] sectored_entries_5_data_0;
  reg [63:0] _RAND_46;
  reg [33:0] sectored_entries_5_data_1;
  reg [63:0] _RAND_47;
  reg [33:0] sectored_entries_5_data_2;
  reg [63:0] _RAND_48;
  reg [33:0] sectored_entries_5_data_3;
  reg [63:0] _RAND_49;
  reg  sectored_entries_5_valid_0;
  reg [31:0] _RAND_50;
  reg  sectored_entries_5_valid_1;
  reg [31:0] _RAND_51;
  reg  sectored_entries_5_valid_2;
  reg [31:0] _RAND_52;
  reg  sectored_entries_5_valid_3;
  reg [31:0] _RAND_53;
  reg [19:0] sectored_entries_6_tag;
  reg [31:0] _RAND_54;
  reg [33:0] sectored_entries_6_data_0;
  reg [63:0] _RAND_55;
  reg [33:0] sectored_entries_6_data_1;
  reg [63:0] _RAND_56;
  reg [33:0] sectored_entries_6_data_2;
  reg [63:0] _RAND_57;
  reg [33:0] sectored_entries_6_data_3;
  reg [63:0] _RAND_58;
  reg  sectored_entries_6_valid_0;
  reg [31:0] _RAND_59;
  reg  sectored_entries_6_valid_1;
  reg [31:0] _RAND_60;
  reg  sectored_entries_6_valid_2;
  reg [31:0] _RAND_61;
  reg  sectored_entries_6_valid_3;
  reg [31:0] _RAND_62;
  reg [19:0] sectored_entries_7_tag;
  reg [31:0] _RAND_63;
  reg [33:0] sectored_entries_7_data_0;
  reg [63:0] _RAND_64;
  reg [33:0] sectored_entries_7_data_1;
  reg [63:0] _RAND_65;
  reg [33:0] sectored_entries_7_data_2;
  reg [63:0] _RAND_66;
  reg [33:0] sectored_entries_7_data_3; 
  reg [63:0] _RAND_67;
  reg  sectored_entries_7_valid_0;
  reg [31:0] _RAND_68;
  reg  sectored_entries_7_valid_1;
  reg [31:0] _RAND_69;
  reg  sectored_entries_7_valid_2;
  reg [31:0] _RAND_70;
  reg  sectored_entries_7_valid_3;
  reg [31:0] _RAND_71;
  reg [19:0] superpage_entries_0_tag;
  reg [31:0] _RAND_72;
  reg [33:0] superpage_entries_0_data_0;
  reg [63:0] _RAND_73;
  reg  superpage_entries_0_valid_0;
  reg [31:0] _RAND_74;
  reg [19:0] superpage_entries_1_tag;
  reg [31:0] _RAND_75;
  reg [33:0] superpage_entries_1_data_0;
  reg [63:0] _RAND_76;
  reg  superpage_entries_1_valid_0;
  reg [31:0] _RAND_77;
  reg [19:0] superpage_entries_2_tag;
  reg [31:0] _RAND_78;
  reg [33:0] superpage_entries_2_data_0;
  reg [63:0] _RAND_79;
  reg  superpage_entries_2_valid_0;
  reg [31:0] _RAND_80;
  reg [19:0] superpage_entries_3_tag;
  reg [31:0] _RAND_81;
  reg [33:0] superpage_entries_3_data_0;
  reg [63:0] _RAND_82;
  reg  superpage_entries_3_valid_0;
  reg [31:0] _RAND_83;
  reg  special_entry_level;
  reg [31:0] _RAND_84;
  reg [19:0] special_entry_tag;
  reg [31:0] _RAND_85;
  reg [33:0] special_entry_data_0;
  reg [63:0] _RAND_86;
  reg  special_entry_valid_0;
  reg [31:0] _RAND_87;
  reg [1:0] state;
  reg [31:0] _RAND_88;
  reg [19:0] r_refill_tag;
  reg [31:0] _RAND_89;
  reg [1:0] r_superpage_repl_addr;
  reg [31:0] _RAND_90;
  reg [2:0] r_sectored_repl_addr;
  reg [31:0] _RAND_91;
  reg [2:0] r_sectored_hit_addr;
  reg [31:0] _RAND_92;
  reg  r_sectored_hit;
  reg [31:0] _RAND_93;
  wire  priv_s;
  wire  priv_uses_vm;
  wire  vm_enabled;
  wire [19:0] vpn;
  wire [19:0] refill_ppn;
  wire  invalidate_refill;
  wire [19:0] mpu_ppn;
  wire [31:0] mpu_physaddr;
  wire [2:0] mpu_priv;
  wire  legal_address;
  wire  cacheable;
  wire  deny_access_to_debug;
  wire  prot_r;
  wire  prot_w;
  wire  prot_al; 
  wire  prot_x;
  wire  prot_eff;
  wire  sector_hits_0;
  wire  sector_hits_1;
  wire  sector_hits_2;
  wire  sector_hits_3;
  wire  sector_hits_4;
  wire  sector_hits_5;
  wire  sector_hits_6; 
  wire  sector_hits_7;
  wire  superpage_hits_0;
  wire  superpage_hits_1;
  wire  superpage_hits_2;
  wire  superpage_hits_3;
  wire  hitsVec_0;
  wire  hitsVec_1;
  wire  hitsVec_2;
  wire  hitsVec_3;
  wire  hitsVec_4;
  wire  hitsVec_5;
  wire  hitsVec_6;
  wire  hitsVec_7;
  wire  hitsVec_8;
  wire  hitsVec_9;
  wire  hitsVec_10;
  wire  hitsVec_11;
  wire  hitsVec_12;
  wire [12:0] real_hits;
  wire [13:0] hits;
  wire [19:0] ppn;
  wire [13:0] ptw_ae_array;
  wire [12:0] priv_rw_ok; 
  wire [13:0] r_array;
  wire [13:0] w_array;
  wire [13:0] pr_array;
  wire [13:0] pw_array;
  wire [13:0] eff_array;
  wire [13:0] c_array;
  wire [13:0] paa_array;
  wire [13:0] pal_array;
  wire [13:0] paa_array_if_cached;
  wire [13:0] pal_array_if_cached;
  wire  misaligned;
  wire  cmd_lrsc;
  wire  cmd_amo_logical;
  wire  cmd_amo_arithmetic;
  wire  cmd_read;
  wire  cmd_write;
  wire  cmd_write_perms;
  wire [13:0] ae_array;
  wire [13:0] ae_ld_array;
  wire [13:0] ae_st_array;
  wire [13:0] ma_ld_array;
  wire [13:0] ma_st_array; 
  wire [13:0] pf_ld_array;
  wire [13:0] pf_st_array;
  wire  tlb_hit;
  wire  tlb_miss;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  wire  multipleHits;
  reg [6:0] _T_1904;
  reg [2:0] _T_1905;
  _2_1 _2 (
    .io_x_ppn(_2_io_x_ppn),
    .io_x_u(_2_io_x_u),
    .io_x_ae(_2_io_x_ae),
    .io_x_sw(_2_io_x_sw),
    .io_x_sx(_2_io_x_sx),
    .io_x_sr(_2_io_x_sr),
    .io_x_pw(_2_io_x_pw),
    .io_x_px(_2_io_x_px),
    .io_x_pr(_2_io_x_pr),
    .io_x_pal(_2_io_x_pal),
    .io_x_paa(_2_io_x_paa),
    .io_x_eff(_2_io_x_eff),
    .io_x_c(_2_io_x_c),
    .io_y_ppn(_2_io_y_ppn),
    .io_y_u(_2_io_y_u),
    .io_y_ae(_2_io_y_ae),
    .io_y_sw(_2_io_y_sw),
    .io_y_sx(_2_io_y_sx),
    .io_y_sr(_2_io_y_sr),
    .io_y_pw(_2_io_y_pw),
    .io_y_px(_2_io_y_px),
    .io_y_pr(_2_io_y_pr),
    .io_y_pal(_2_io_y_pal),
    .io_y_paa(_2_io_y_paa),
    .io_y_eff(_2_io_y_eff),
    .io_y_c(_2_io_y_c)
  );
  PMPChecker pmp (
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x)
  );
  _2_1 _2_1 ( 
    .io_x_ppn(_2_1_io_x_ppn),
    .io_x_u(_2_1_io_x_u),
    .io_x_ae(_2_1_io_x_ae),
    .io_x_sw(_2_1_io_x_sw),
    .io_x_sx(_2_1_io_x_sx),
    .io_x_sr(_2_1_io_x_sr),
    .io_x_pw(_2_1_io_x_pw),
    .io_x_px(_2_1_io_x_px),
    .io_x_pr(_2_1_io_x_pr),
    .io_x_pal(_2_1_io_x_pal),
    .io_x_paa(_2_1_io_x_paa),
    .io_x_eff(_2_1_io_x_eff),
    .io_x_c(_2_1_io_x_c),
    .io_y_ppn(_2_1_io_y_ppn),
    .io_y_u(_2_1_io_y_u),
    .io_y_ae(_2_1_io_y_ae),
    .io_y_sw(_2_1_io_y_sw),
    .io_y_sx(_2_1_io_y_sx),
    .io_y_sr(_2_1_io_y_sr),
    .io_y_pw(_2_1_io_y_pw),
    .io_y_px(_2_1_io_y_px),
    .io_y_pr(_2_1_io_y_pr),
    .io_y_pal(_2_1_io_y_pal),
    .io_y_paa(_2_1_io_y_paa),
    .io_y_eff(_2_1_io_y_eff),
    .io_y_c(_2_1_io_y_c)
  );
  _2_1 _2_2 (
    .io_x_ppn(_2_2_io_x_ppn),
    .io_x_u(_2_2_io_x_u),
    .io_x_ae(_2_2_io_x_ae),
    .io_x_sw(_2_2_io_x_sw),
    .io_x_sx(_2_2_io_x_sx),
    .io_x_sr(_2_2_io_x_sr),
    .io_x_pw(_2_2_io_x_pw),
    .io_x_px(_2_2_io_x_px),
    .io_x_pr(_2_2_io_x_pr),
    .io_x_pal(_2_2_io_x_pal),
    .io_x_paa(_2_2_io_x_paa),
    .io_x_eff(_2_2_io_x_eff),
    .io_x_c(_2_2_io_x_c),
    .io_y_ppn(_2_2_io_y_ppn),
    .io_y_u(_2_2_io_y_u),
    .io_y_ae(_2_2_io_y_ae),
    .io_y_sw(_2_2_io_y_sw),
    .io_y_sx(_2_2_io_y_sx),
    .io_y_sr(_2_2_io_y_sr),
    .io_y_pw(_2_2_io_y_pw),
    .io_y_px(_2_2_io_y_px),
    .io_y_pr(_2_2_io_y_pr),
    .io_y_pal(_2_2_io_y_pal),
    .io_y_paa(_2_2_io_y_paa),
    .io_y_eff(_2_2_io_y_eff),
    .io_y_c(_2_2_io_y_c)
  );
  _2_1 _2_3 (
    .io_x_ppn(_2_3_io_x_ppn),
    .io_x_u(_2_3_io_x_u),
    .io_x_ae(_2_3_io_x_ae),
    .io_x_sw(_2_3_io_x_sw),
    .io_x_sx(_2_3_io_x_sx),
    .io_x_sr(_2_3_io_x_sr),
    .io_x_pw(_2_3_io_x_pw),
    .io_x_px(_2_3_io_x_px),
    .io_x_pr(_2_3_io_x_pr),
    .io_x_pal(_2_3_io_x_pal),
    .io_x_paa(_2_3_io_x_paa),
    .io_x_eff(_2_3_io_x_eff),
    .io_x_c(_2_3_io_x_c),
    .io_y_ppn(_2_3_io_y_ppn),
    .io_y_u(_2_3_io_y_u),
    .io_y_ae(_2_3_io_y_ae),
    .io_y_sw(_2_3_io_y_sw),
    .io_y_sx(_2_3_io_y_sx),
    .io_y_sr(_2_3_io_y_sr),
    .io_y_pw(_2_3_io_y_pw),
    .io_y_px(_2_3_io_y_px),
    .io_y_pr(_2_3_io_y_pr),
    .io_y_pal(_2_3_io_y_pal),
    .io_y_paa(_2_3_io_y_paa),
    .io_y_eff(_2_3_io_y_eff),
    .io_y_c(_2_3_io_y_c)
  );
  _2_1 _2_4 (
    .io_x_ppn(_2_4_io_x_ppn),
    .io_x_u(_2_4_io_x_u),
    .io_x_ae(_2_4_io_x_ae),
    .io_x_sw(_2_4_io_x_sw),
    .io_x_sx(_2_4_io_x_sx),
    .io_x_sr(_2_4_io_x_sr),
    .io_x_pw(_2_4_io_x_pw),
    .io_x_px(_2_4_io_x_px),
    .io_x_pr(_2_4_io_x_pr),
    .io_x_pal(_2_4_io_x_pal),
    .io_x_paa(_2_4_io_x_paa),
    .io_x_eff(_2_4_io_x_eff),
    .io_x_c(_2_4_io_x_c),
    .io_y_ppn(_2_4_io_y_ppn),
    .io_y_u(_2_4_io_y_u),
    .io_y_ae(_2_4_io_y_ae),
    .io_y_sw(_2_4_io_y_sw),
    .io_y_sx(_2_4_io_y_sx),
    .io_y_sr(_2_4_io_y_sr),
    .io_y_pw(_2_4_io_y_pw),
    .io_y_px(_2_4_io_y_px),
    .io_y_pr(_2_4_io_y_pr),
    .io_y_pal(_2_4_io_y_pal),
    .io_y_paa(_2_4_io_y_paa),
    .io_y_eff(_2_4_io_y_eff),
    .io_y_c(_2_4_io_y_c)
  );
  _2_1 _2_5 ( 
    .io_x_ppn(_2_5_io_x_ppn),
    .io_x_u(_2_5_io_x_u),
    .io_x_ae(_2_5_io_x_ae),
    .io_x_sw(_2_5_io_x_sw),
    .io_x_sx(_2_5_io_x_sx),
    .io_x_sr(_2_5_io_x_sr),
    .io_x_pw(_2_5_io_x_pw),
    .io_x_px(_2_5_io_x_px),
    .io_x_pr(_2_5_io_x_pr),
    .io_x_pal(_2_5_io_x_pal),
    .io_x_paa(_2_5_io_x_paa),
    .io_x_eff(_2_5_io_x_eff),
    .io_x_c(_2_5_io_x_c),
    .io_y_ppn(_2_5_io_y_ppn),
    .io_y_u(_2_5_io_y_u),
    .io_y_ae(_2_5_io_y_ae),
    .io_y_sw(_2_5_io_y_sw),
    .io_y_sx(_2_5_io_y_sx),
    .io_y_sr(_2_5_io_y_sr),
    .io_y_pw(_2_5_io_y_pw),
    .io_y_px(_2_5_io_y_px),
    .io_y_pr(_2_5_io_y_pr),
    .io_y_pal(_2_5_io_y_pal),
    .io_y_paa(_2_5_io_y_paa),
    .io_y_eff(_2_5_io_y_eff),
    .io_y_c(_2_5_io_y_c)
  );
  _2_1 _2_6 (
    .io_x_ppn(_2_6_io_x_ppn),
    .io_x_u(_2_6_io_x_u),
    .io_x_ae(_2_6_io_x_ae),
    .io_x_sw(_2_6_io_x_sw),
    .io_x_sx(_2_6_io_x_sx),
    .io_x_sr(_2_6_io_x_sr),
    .io_x_pw(_2_6_io_x_pw),
    .io_x_px(_2_6_io_x_px),
    .io_x_pr(_2_6_io_x_pr),
    .io_x_pal(_2_6_io_x_pal),
    .io_x_paa(_2_6_io_x_paa),
    .io_x_eff(_2_6_io_x_eff),
    .io_x_c(_2_6_io_x_c),
    .io_y_ppn(_2_6_io_y_ppn),
    .io_y_u(_2_6_io_y_u),
    .io_y_ae(_2_6_io_y_ae),
    .io_y_sw(_2_6_io_y_sw),
    .io_y_sx(_2_6_io_y_sx),
    .io_y_sr(_2_6_io_y_sr),
    .io_y_pw(_2_6_io_y_pw),
    .io_y_px(_2_6_io_y_px),
    .io_y_pr(_2_6_io_y_pr),
    .io_y_pal(_2_6_io_y_pal),
    .io_y_paa(_2_6_io_y_paa),
    .io_y_eff(_2_6_io_y_eff),
    .io_y_c(_2_6_io_y_c)
  );
  _2_1 _2_7 (
    .io_x_ppn(_2_7_io_x_ppn),
    .io_x_u(_2_7_io_x_u),
    .io_x_ae(_2_7_io_x_ae),
    .io_x_sw(_2_7_io_x_sw),
    .io_x_sx(_2_7_io_x_sx),
    .io_x_sr(_2_7_io_x_sr),
    .io_x_pw(_2_7_io_x_pw),
    .io_x_px(_2_7_io_x_px),
    .io_x_pr(_2_7_io_x_pr),
    .io_x_pal(_2_7_io_x_pal),
    .io_x_paa(_2_7_io_x_paa),
    .io_x_eff(_2_7_io_x_eff),
    .io_x_c(_2_7_io_x_c),
    .io_y_ppn(_2_7_io_y_ppn),
    .io_y_u(_2_7_io_y_u),
    .io_y_ae(_2_7_io_y_ae),
    .io_y_sw(_2_7_io_y_sw),
    .io_y_sx(_2_7_io_y_sx),
    .io_y_sr(_2_7_io_y_sr),
    .io_y_pw(_2_7_io_y_pw),
    .io_y_px(_2_7_io_y_px),
    .io_y_pr(_2_7_io_y_pr),
    .io_y_pal(_2_7_io_y_pal),
    .io_y_paa(_2_7_io_y_paa),
    .io_y_eff(_2_7_io_y_eff),
    .io_y_c(_2_7_io_y_c)
  );
  _2_1 _2_8 (
    .io_x_ppn(_2_8_io_x_ppn),
    .io_x_u(_2_8_io_x_u),
    .io_x_ae(_2_8_io_x_ae),
    .io_x_sw(_2_8_io_x_sw),
    .io_x_sx(_2_8_io_x_sx),
    .io_x_sr(_2_8_io_x_sr),
    .io_x_pw(_2_8_io_x_pw),
    .io_x_px(_2_8_io_x_px),
    .io_x_pr(_2_8_io_x_pr),
    .io_x_pal(_2_8_io_x_pal),
    .io_x_paa(_2_8_io_x_paa),
    .io_x_eff(_2_8_io_x_eff),
    .io_x_c(_2_8_io_x_c),
    .io_y_ppn(_2_8_io_y_ppn),
    .io_y_u(_2_8_io_y_u),
    .io_y_ae(_2_8_io_y_ae),
    .io_y_sw(_2_8_io_y_sw),
    .io_y_sx(_2_8_io_y_sx),
    .io_y_sr(_2_8_io_y_sr),
    .io_y_pw(_2_8_io_y_pw),
    .io_y_px(_2_8_io_y_px),
    .io_y_pr(_2_8_io_y_pr),
    .io_y_pal(_2_8_io_y_pal),
    .io_y_paa(_2_8_io_y_paa),
    .io_y_eff(_2_8_io_y_eff),
    .io_y_c(_2_8_io_y_c)
  );
  _2_1 _2_9 (
    .io_x_ppn(_2_9_io_x_ppn),
    .io_x_u(_2_9_io_x_u),
    .io_x_ae(_2_9_io_x_ae),
    .io_x_sw(_2_9_io_x_sw),
    .io_x_sx(_2_9_io_x_sx),
    .io_x_sr(_2_9_io_x_sr),
    .io_x_pw(_2_9_io_x_pw),
    .io_x_px(_2_9_io_x_px),
    .io_x_pr(_2_9_io_x_pr),
    .io_x_pal(_2_9_io_x_pal),
    .io_x_paa(_2_9_io_x_paa),
    .io_x_eff(_2_9_io_x_eff),
    .io_x_c(_2_9_io_x_c),
    .io_y_ppn(_2_9_io_y_ppn),
    .io_y_u(_2_9_io_y_u),
    .io_y_ae(_2_9_io_y_ae),
    .io_y_sw(_2_9_io_y_sw),
    .io_y_sx(_2_9_io_y_sx),
    .io_y_sr(_2_9_io_y_sr),
    .io_y_pw(_2_9_io_y_pw),
    .io_y_px(_2_9_io_y_px),
    .io_y_pr(_2_9_io_y_pr),
    .io_y_pal(_2_9_io_y_pal),
    .io_y_paa(_2_9_io_y_paa),
    .io_y_eff(_2_9_io_y_eff),
    .io_y_c(_2_9_io_y_c)
  );
  _2_1 _2_10 (
    .io_x_ppn(_2_10_io_x_ppn),
    .io_x_u(_2_10_io_x_u),
    .io_x_ae(_2_10_io_x_ae),
    .io_x_sw(_2_10_io_x_sw),
    .io_x_sx(_2_10_io_x_sx),
    .io_x_sr(_2_10_io_x_sr),
    .io_x_pw(_2_10_io_x_pw),
    .io_x_px(_2_10_io_x_px),
    .io_x_pr(_2_10_io_x_pr),
    .io_x_pal(_2_10_io_x_pal),
    .io_x_paa(_2_10_io_x_paa),
    .io_x_eff(_2_10_io_x_eff),
    .io_x_c(_2_10_io_x_c),
    .io_y_ppn(_2_10_io_y_ppn),
    .io_y_u(_2_10_io_y_u),
    .io_y_ae(_2_10_io_y_ae),
    .io_y_sw(_2_10_io_y_sw),
    .io_y_sx(_2_10_io_y_sx),
    .io_y_sr(_2_10_io_y_sr),
    .io_y_pw(_2_10_io_y_pw),
    .io_y_px(_2_10_io_y_px),
    .io_y_pr(_2_10_io_y_pr),
    .io_y_pal(_2_10_io_y_pal),
    .io_y_paa(_2_10_io_y_paa),
    .io_y_eff(_2_10_io_y_eff),
    .io_y_c(_2_10_io_y_c)
  );
  _2_1 _2_11 (
    .io_x_ppn(_2_11_io_x_ppn),
    .io_x_u(_2_11_io_x_u),
    .io_x_ae(_2_11_io_x_ae),
    .io_x_sw(_2_11_io_x_sw),
    .io_x_sx(_2_11_io_x_sx),
    .io_x_sr(_2_11_io_x_sr),
    .io_x_pw(_2_11_io_x_pw),
    .io_x_px(_2_11_io_x_px),
    .io_x_pr(_2_11_io_x_pr),
    .io_x_pal(_2_11_io_x_pal),
    .io_x_paa(_2_11_io_x_paa),
    .io_x_eff(_2_11_io_x_eff),
    .io_x_c(_2_11_io_x_c),
    .io_y_ppn(_2_11_io_y_ppn),
    .io_y_u(_2_11_io_y_u),
    .io_y_ae(_2_11_io_y_ae),
    .io_y_sw(_2_11_io_y_sw),
    .io_y_sx(_2_11_io_y_sx),
    .io_y_sr(_2_11_io_y_sr),
    .io_y_pw(_2_11_io_y_pw),
    .io_y_px(_2_11_io_y_px),
    .io_y_pr(_2_11_io_y_pr),
    .io_y_pal(_2_11_io_y_pal),
    .io_y_paa(_2_11_io_y_paa),
    .io_y_eff(_2_11_io_y_eff),
    .io_y_c(_2_11_io_y_c)
  );
  _2_1 _2_12 (
    .io_x_ppn(_2_12_io_x_ppn),
    .io_x_u(_2_12_io_x_u),
    .io_x_ae(_2_12_io_x_ae),
    .io_x_sw(_2_12_io_x_sw),
    .io_x_sx(_2_12_io_x_sx),
    .io_x_sr(_2_12_io_x_sr),
    .io_x_pw(_2_12_io_x_pw),
    .io_x_px(_2_12_io_x_px),
    .io_x_pr(_2_12_io_x_pr),
    .io_x_pal(_2_12_io_x_pal),
    .io_x_paa(_2_12_io_x_paa),
    .io_x_eff(_2_12_io_x_eff),
    .io_x_c(_2_12_io_x_c),
    .io_y_ppn(_2_12_io_y_ppn),
    .io_y_u(_2_12_io_y_u),
    .io_y_ae(_2_12_io_y_ae),
    .io_y_sw(_2_12_io_y_sw),
    .io_y_sx(_2_12_io_y_sx),
    .io_y_sr(_2_12_io_y_sr),
    .io_y_pw(_2_12_io_y_pw),
    .io_y_px(_2_12_io_y_px),
    .io_y_pr(_2_12_io_y_pr),
    .io_y_pal(_2_12_io_y_pal),
    .io_y_paa(_2_12_io_y_paa),
    .io_y_eff(_2_12_io_y_eff),
    .io_y_c(_2_12_io_y_c)
  );
  _2_1 _2_13 (
    .io_x_ppn(_2_13_io_x_ppn),
    .io_x_u(_2_13_io_x_u),
    .io_x_ae(_2_13_io_x_ae),
    .io_x_sw(_2_13_io_x_sw),
    .io_x_sx(_2_13_io_x_sx),
    .io_x_sr(_2_13_io_x_sr),
    .io_x_pw(_2_13_io_x_pw),
    .io_x_px(_2_13_io_x_px),
    .io_x_pr(_2_13_io_x_pr),
    .io_x_pal(_2_13_io_x_pal),
    .io_x_paa(_2_13_io_x_paa),
    .io_x_eff(_2_13_io_x_eff),
    .io_x_c(_2_13_io_x_c),
    .io_y_ppn(_2_13_io_y_ppn),
    .io_y_u(_2_13_io_y_u),
    .io_y_ae(_2_13_io_y_ae),
    .io_y_sw(_2_13_io_y_sw),
    .io_y_sx(_2_13_io_y_sx),
    .io_y_sr(_2_13_io_y_sr),
    .io_y_pw(_2_13_io_y_pw),
    .io_y_px(_2_13_io_y_px),
    .io_y_pr(_2_13_io_y_pr),
    .io_y_pal(_2_13_io_y_pal),
    .io_y_paa(_2_13_io_y_paa),
    .io_y_eff(_2_13_io_y_eff),
    .io_y_c(_2_13_io_y_c)
  );
  _2_1 _2_14 (
    .io_x_ppn(_2_14_io_x_ppn),
    .io_x_u(_2_14_io_x_u),
    .io_x_ae(_2_14_io_x_ae),
    .io_x_sw(_2_14_io_x_sw),
    .io_x_sx(_2_14_io_x_sx),
    .io_x_sr(_2_14_io_x_sr),
    .io_x_pw(_2_14_io_x_pw),
    .io_x_px(_2_14_io_x_px),
    .io_x_pr(_2_14_io_x_pr),
    .io_x_pal(_2_14_io_x_pal),
    .io_x_paa(_2_14_io_x_paa),
    .io_x_eff(_2_14_io_x_eff),
    .io_x_c(_2_14_io_x_c),
    .io_y_ppn(_2_14_io_y_ppn),
    .io_y_u(_2_14_io_y_u),
    .io_y_ae(_2_14_io_y_ae),
    .io_y_sw(_2_14_io_y_sw),
    .io_y_sx(_2_14_io_y_sx),
    .io_y_sr(_2_14_io_y_sr),
    .io_y_pw(_2_14_io_y_pw),
    .io_y_px(_2_14_io_y_px),
    .io_y_pr(_2_14_io_y_pr),
    .io_y_pal(_2_14_io_y_pal),
    .io_y_paa(_2_14_io_y_paa),
    .io_y_eff(_2_14_io_y_eff),
    .io_y_c(_2_14_io_y_c)
  );
  _2_1 _2_15 (
    .io_x_ppn(_2_15_io_x_ppn),
    .io_x_u(_2_15_io_x_u),
    .io_x_ae(_2_15_io_x_ae),
    .io_x_sw(_2_15_io_x_sw),
    .io_x_sx(_2_15_io_x_sx),
    .io_x_sr(_2_15_io_x_sr),
    .io_x_pw(_2_15_io_x_pw),
    .io_x_px(_2_15_io_x_px),
    .io_x_pr(_2_15_io_x_pr),
    .io_x_pal(_2_15_io_x_pal),
    .io_x_paa(_2_15_io_x_paa),
    .io_x_eff(_2_15_io_x_eff),
    .io_x_c(_2_15_io_x_c),
    .io_y_ppn(_2_15_io_y_ppn),
    .io_y_u(_2_15_io_y_u),
    .io_y_ae(_2_15_io_y_ae),
    .io_y_sw(_2_15_io_y_sw),
    .io_y_sx(_2_15_io_y_sx),
    .io_y_sr(_2_15_io_y_sr),
    .io_y_pw(_2_15_io_y_pw),
    .io_y_px(_2_15_io_y_px),
    .io_y_pr(_2_15_io_y_pr),
    .io_y_pal(_2_15_io_y_pal),
    .io_y_paa(_2_15_io_y_paa),
    .io_y_eff(_2_15_io_y_eff),
    .io_y_c(_2_15_io_y_c)
  );
  _2_1 _2_16 (
    .io_x_ppn(_2_16_io_x_ppn),
    .io_x_u(_2_16_io_x_u),
    .io_x_ae(_2_16_io_x_ae),
    .io_x_sw(_2_16_io_x_sw),
    .io_x_sx(_2_16_io_x_sx),
    .io_x_sr(_2_16_io_x_sr),
    .io_x_pw(_2_16_io_x_pw),
    .io_x_px(_2_16_io_x_px),
    .io_x_pr(_2_16_io_x_pr),
    .io_x_pal(_2_16_io_x_pal),
    .io_x_paa(_2_16_io_x_paa),
    .io_x_eff(_2_16_io_x_eff),
    .io_x_c(_2_16_io_x_c),
    .io_y_ppn(_2_16_io_y_ppn),
    .io_y_u(_2_16_io_y_u),
    .io_y_ae(_2_16_io_y_ae),
    .io_y_sw(_2_16_io_y_sw),
    .io_y_sx(_2_16_io_y_sx),
    .io_y_sr(_2_16_io_y_sr),
    .io_y_pw(_2_16_io_y_pw),
    .io_y_px(_2_16_io_y_px),
    .io_y_pr(_2_16_io_y_pr),
    .io_y_pal(_2_16_io_y_pal),
    .io_y_paa(_2_16_io_y_paa),
    .io_y_eff(_2_16_io_y_eff),
    .io_y_c(_2_16_io_y_c)
  );
  _2_1 _2_17 ( 
    .io_x_ppn(_2_17_io_x_ppn),
    .io_x_u(_2_17_io_x_u),
    .io_x_ae(_2_17_io_x_ae),
    .io_x_sw(_2_17_io_x_sw),
    .io_x_sx(_2_17_io_x_sx),
    .io_x_sr(_2_17_io_x_sr),
    .io_x_pw(_2_17_io_x_pw),
    .io_x_px(_2_17_io_x_px),
    .io_x_pr(_2_17_io_x_pr),
    .io_x_pal(_2_17_io_x_pal),
    .io_x_paa(_2_17_io_x_paa),
    .io_x_eff(_2_17_io_x_eff),
    .io_x_c(_2_17_io_x_c),
    .io_y_ppn(_2_17_io_y_ppn),
    .io_y_u(_2_17_io_y_u),
    .io_y_ae(_2_17_io_y_ae),
    .io_y_sw(_2_17_io_y_sw),
    .io_y_sx(_2_17_io_y_sx),
    .io_y_sr(_2_17_io_y_sr),
    .io_y_pw(_2_17_io_y_pw),
    .io_y_px(_2_17_io_y_px),
    .io_y_pr(_2_17_io_y_pr),
    .io_y_pal(_2_17_io_y_pal),
    .io_y_paa(_2_17_io_y_paa),
    .io_y_eff(_2_17_io_y_eff),
    .io_y_c(_2_17_io_y_c)
  );
  _2_1 _2_18 (
    .io_x_ppn(_2_18_io_x_ppn),
    .io_x_u(_2_18_io_x_u),
    .io_x_ae(_2_18_io_x_ae),
    .io_x_sw(_2_18_io_x_sw),
    .io_x_sx(_2_18_io_x_sx),
    .io_x_sr(_2_18_io_x_sr),
    .io_x_pw(_2_18_io_x_pw),
    .io_x_px(_2_18_io_x_px),
    .io_x_pr(_2_18_io_x_pr),
    .io_x_pal(_2_18_io_x_pal),
    .io_x_paa(_2_18_io_x_paa),
    .io_x_eff(_2_18_io_x_eff),
    .io_x_c(_2_18_io_x_c),
    .io_y_ppn(_2_18_io_y_ppn),
    .io_y_u(_2_18_io_y_u),
    .io_y_ae(_2_18_io_y_ae),
    .io_y_sw(_2_18_io_y_sw),
    .io_y_sx(_2_18_io_y_sx),
    .io_y_sr(_2_18_io_y_sr),
    .io_y_pw(_2_18_io_y_pw),
    .io_y_px(_2_18_io_y_px),
    .io_y_pr(_2_18_io_y_pr),
    .io_y_pal(_2_18_io_y_pal),
    .io_y_paa(_2_18_io_y_paa),
    .io_y_eff(_2_18_io_y_eff),
    .io_y_c(_2_18_io_y_c)
  );
  _2_1 _2_19 (
    .io_x_ppn(_2_19_io_x_ppn),
    .io_x_u(_2_19_io_x_u),
    .io_x_ae(_2_19_io_x_ae),
    .io_x_sw(_2_19_io_x_sw),
    .io_x_sx(_2_19_io_x_sx),
    .io_x_sr(_2_19_io_x_sr),
    .io_x_pw(_2_19_io_x_pw),
    .io_x_px(_2_19_io_x_px),
    .io_x_pr(_2_19_io_x_pr),
    .io_x_pal(_2_19_io_x_pal),
    .io_x_paa(_2_19_io_x_paa),
    .io_x_eff(_2_19_io_x_eff),
    .io_x_c(_2_19_io_x_c),
    .io_y_ppn(_2_19_io_y_ppn),
    .io_y_u(_2_19_io_y_u),
    .io_y_ae(_2_19_io_y_ae),
    .io_y_sw(_2_19_io_y_sw),
    .io_y_sx(_2_19_io_y_sx),
    .io_y_sr(_2_19_io_y_sr),
    .io_y_pw(_2_19_io_y_pw),
    .io_y_px(_2_19_io_y_px),
    .io_y_pr(_2_19_io_y_pr),
    .io_y_pal(_2_19_io_y_pal),
    .io_y_paa(_2_19_io_y_paa),
    .io_y_eff(_2_19_io_y_eff),
    .io_y_c(_2_19_io_y_c)
  );
  _2_1 _2_20 (
    .io_x_ppn(_2_20_io_x_ppn),
    .io_x_u(_2_20_io_x_u),
    .io_x_ae(_2_20_io_x_ae),
    .io_x_sw(_2_20_io_x_sw),
    .io_x_sx(_2_20_io_x_sx),
    .io_x_sr(_2_20_io_x_sr),
    .io_x_pw(_2_20_io_x_pw),
    .io_x_px(_2_20_io_x_px),
    .io_x_pr(_2_20_io_x_pr),
    .io_x_pal(_2_20_io_x_pal),
    .io_x_paa(_2_20_io_x_paa),
    .io_x_eff(_2_20_io_x_eff),
    .io_x_c(_2_20_io_x_c),
    .io_y_ppn(_2_20_io_y_ppn),
    .io_y_u(_2_20_io_y_u),
    .io_y_ae(_2_20_io_y_ae),
    .io_y_sw(_2_20_io_y_sw),
    .io_y_sx(_2_20_io_y_sx),
    .io_y_sr(_2_20_io_y_sr),
    .io_y_pw(_2_20_io_y_pw),
    .io_y_px(_2_20_io_y_px),
    .io_y_pr(_2_20_io_y_pr),
    .io_y_pal(_2_20_io_y_pal),
    .io_y_paa(_2_20_io_y_paa),
    .io_y_eff(_2_20_io_y_eff),
    .io_y_c(_2_20_io_y_c)
  );
  _2_1 _2_21 (
    .io_x_ppn(_2_21_io_x_ppn),
    .io_x_u(_2_21_io_x_u),
    .io_x_ae(_2_21_io_x_ae),
    .io_x_sw(_2_21_io_x_sw),
    .io_x_sx(_2_21_io_x_sx),
    .io_x_sr(_2_21_io_x_sr),
    .io_x_pw(_2_21_io_x_pw),
    .io_x_px(_2_21_io_x_px),
    .io_x_pr(_2_21_io_x_pr),
    .io_x_pal(_2_21_io_x_pal),
    .io_x_paa(_2_21_io_x_paa),
    .io_x_eff(_2_21_io_x_eff),
    .io_x_c(_2_21_io_x_c),
    .io_y_ppn(_2_21_io_y_ppn),
    .io_y_u(_2_21_io_y_u),
    .io_y_ae(_2_21_io_y_ae),
    .io_y_sw(_2_21_io_y_sw),
    .io_y_sx(_2_21_io_y_sx),
    .io_y_sr(_2_21_io_y_sr),
    .io_y_pw(_2_21_io_y_pw),
    .io_y_px(_2_21_io_y_px),
    .io_y_pr(_2_21_io_y_pr),
    .io_y_pal(_2_21_io_y_pal),
    .io_y_paa(_2_21_io_y_paa),
    .io_y_eff(_2_21_io_y_eff),
    .io_y_c(_2_21_io_y_c)
  );
  _2_1 _2_22 (
    .io_x_ppn(_2_22_io_x_ppn),
    .io_x_u(_2_22_io_x_u),
    .io_x_ae(_2_22_io_x_ae),
    .io_x_sw(_2_22_io_x_sw),
    .io_x_sx(_2_22_io_x_sx),
    .io_x_sr(_2_22_io_x_sr),
    .io_x_pw(_2_22_io_x_pw),
    .io_x_px(_2_22_io_x_px),
    .io_x_pr(_2_22_io_x_pr),
    .io_x_pal(_2_22_io_x_pal),
    .io_x_paa(_2_22_io_x_paa),
    .io_x_eff(_2_22_io_x_eff),
    .io_x_c(_2_22_io_x_c),
    .io_y_ppn(_2_22_io_y_ppn),
    .io_y_u(_2_22_io_y_u),
    .io_y_ae(_2_22_io_y_ae),
    .io_y_sw(_2_22_io_y_sw),
    .io_y_sx(_2_22_io_y_sx),
    .io_y_sr(_2_22_io_y_sr),
    .io_y_pw(_2_22_io_y_pw),
    .io_y_px(_2_22_io_y_px),
    .io_y_pr(_2_22_io_y_pr),
    .io_y_pal(_2_22_io_y_pal),
    .io_y_paa(_2_22_io_y_paa),
    .io_y_eff(_2_22_io_y_eff),
    .io_y_c(_2_22_io_y_c)
  );
  _2_1 _2_23 (
    .io_x_ppn(_2_23_io_x_ppn),
    .io_x_u(_2_23_io_x_u),
    .io_x_ae(_2_23_io_x_ae),
    .io_x_sw(_2_23_io_x_sw),
    .io_x_sx(_2_23_io_x_sx),
    .io_x_sr(_2_23_io_x_sr),
    .io_x_pw(_2_23_io_x_pw),
    .io_x_px(_2_23_io_x_px),
    .io_x_pr(_2_23_io_x_pr),
    .io_x_pal(_2_23_io_x_pal),
    .io_x_paa(_2_23_io_x_paa),
    .io_x_eff(_2_23_io_x_eff),
    .io_x_c(_2_23_io_x_c),
    .io_y_ppn(_2_23_io_y_ppn),
    .io_y_u(_2_23_io_y_u),
    .io_y_ae(_2_23_io_y_ae),
    .io_y_sw(_2_23_io_y_sw),
    .io_y_sx(_2_23_io_y_sx),
    .io_y_sr(_2_23_io_y_sr),
    .io_y_pw(_2_23_io_y_pw),
    .io_y_px(_2_23_io_y_px),
    .io_y_pr(_2_23_io_y_pr),
    .io_y_pal(_2_23_io_y_pal),
    .io_y_paa(_2_23_io_y_paa),
    .io_y_eff(_2_23_io_y_eff),
    .io_y_c(_2_23_io_y_c)
  );
  _2_1 _2_24 (
    .io_x_ppn(_2_24_io_x_ppn),
    .io_x_u(_2_24_io_x_u),
    .io_x_ae(_2_24_io_x_ae),
    .io_x_sw(_2_24_io_x_sw),
    .io_x_sx(_2_24_io_x_sx),
    .io_x_sr(_2_24_io_x_sr),
    .io_x_pw(_2_24_io_x_pw),
    .io_x_px(_2_24_io_x_px),
    .io_x_pr(_2_24_io_x_pr),
    .io_x_pal(_2_24_io_x_pal),
    .io_x_paa(_2_24_io_x_paa),
    .io_x_eff(_2_24_io_x_eff),
    .io_x_c(_2_24_io_x_c),
    .io_y_ppn(_2_24_io_y_ppn),
    .io_y_u(_2_24_io_y_u),
    .io_y_ae(_2_24_io_y_ae),
    .io_y_sw(_2_24_io_y_sw),
    .io_y_sx(_2_24_io_y_sx),
    .io_y_sr(_2_24_io_y_sr),
    .io_y_pw(_2_24_io_y_pw),
    .io_y_px(_2_24_io_y_px),
    .io_y_pr(_2_24_io_y_pr),
    .io_y_pal(_2_24_io_y_pal),
    .io_y_paa(_2_24_io_y_paa),
    .io_y_eff(_2_24_io_y_eff),
    .io_y_c(_2_24_io_y_c)
  );
  _2_1 _2_25 (
    .io_x_ppn(_2_25_io_x_ppn),
    .io_x_u(_2_25_io_x_u),
    .io_x_ae(_2_25_io_x_ae),
    .io_x_sw(_2_25_io_x_sw),
    .io_x_sx(_2_25_io_x_sx),
    .io_x_sr(_2_25_io_x_sr),
    .io_x_pw(_2_25_io_x_pw),
    .io_x_px(_2_25_io_x_px),
    .io_x_pr(_2_25_io_x_pr),
    .io_x_pal(_2_25_io_x_pal),
    .io_x_paa(_2_25_io_x_paa),
    .io_x_eff(_2_25_io_x_eff),
    .io_x_c(_2_25_io_x_c),
    .io_y_ppn(_2_25_io_y_ppn),
    .io_y_u(_2_25_io_y_u),
    .io_y_ae(_2_25_io_y_ae),
    .io_y_sw(_2_25_io_y_sw),
    .io_y_sx(_2_25_io_y_sx),
    .io_y_sr(_2_25_io_y_sr),
    .io_y_pw(_2_25_io_y_pw),
    .io_y_px(_2_25_io_y_px),
    .io_y_pr(_2_25_io_y_pr),
    .io_y_pal(_2_25_io_y_pal),
    .io_y_paa(_2_25_io_y_paa),
    .io_y_eff(_2_25_io_y_eff),
    .io_y_c(_2_25_io_y_c)
  );
  _2_1 _2_26 (
    .io_x_ppn(_2_26_io_x_ppn),
    .io_x_u(_2_26_io_x_u),
    .io_x_ae(_2_26_io_x_ae),
    .io_x_sw(_2_26_io_x_sw),
    .io_x_sx(_2_26_io_x_sx),
    .io_x_sr(_2_26_io_x_sr),
    .io_x_pw(_2_26_io_x_pw),
    .io_x_px(_2_26_io_x_px),
    .io_x_pr(_2_26_io_x_pr),
    .io_x_pal(_2_26_io_x_pal),
    .io_x_paa(_2_26_io_x_paa),
    .io_x_eff(_2_26_io_x_eff),
    .io_x_c(_2_26_io_x_c),
    .io_y_ppn(_2_26_io_y_ppn),
    .io_y_u(_2_26_io_y_u),
    .io_y_ae(_2_26_io_y_ae),
    .io_y_sw(_2_26_io_y_sw),
    .io_y_sx(_2_26_io_y_sx),
    .io_y_sr(_2_26_io_y_sr),
    .io_y_pw(_2_26_io_y_pw),
    .io_y_px(_2_26_io_y_px),
    .io_y_pr(_2_26_io_y_pr),
    .io_y_pal(_2_26_io_y_pal),
    .io_y_paa(_2_26_io_y_paa),
    .io_y_eff(_2_26_io_y_eff),
    .io_y_c(_2_26_io_y_c)
  );
  _2_1 _2_27 (
    .io_x_ppn(_2_27_io_x_ppn),
    .io_x_u(_2_27_io_x_u),
    .io_x_ae(_2_27_io_x_ae),
    .io_x_sw(_2_27_io_x_sw),
    .io_x_sx(_2_27_io_x_sx),
    .io_x_sr(_2_27_io_x_sr),
    .io_x_pw(_2_27_io_x_pw),
    .io_x_px(_2_27_io_x_px),
    .io_x_pr(_2_27_io_x_pr),
    .io_x_pal(_2_27_io_x_pal),
    .io_x_paa(_2_27_io_x_paa),
    .io_x_eff(_2_27_io_x_eff),
    .io_x_c(_2_27_io_x_c),
    .io_y_ppn(_2_27_io_y_ppn),
    .io_y_u(_2_27_io_y_u),
    .io_y_ae(_2_27_io_y_ae),
    .io_y_sw(_2_27_io_y_sw),
    .io_y_sx(_2_27_io_y_sx),
    .io_y_sr(_2_27_io_y_sr),
    .io_y_pw(_2_27_io_y_pw),
    .io_y_px(_2_27_io_y_px),
    .io_y_pr(_2_27_io_y_pr),
    .io_y_pal(_2_27_io_y_pal),
    .io_y_paa(_2_27_io_y_paa),
    .io_y_eff(_2_27_io_y_eff),
    .io_y_c(_2_27_io_y_c)
  );
  _2_1 _2_28 (
    .io_x_ppn(_2_28_io_x_ppn),
    .io_x_u(_2_28_io_x_u),
    .io_x_ae(_2_28_io_x_ae),
    .io_x_sw(_2_28_io_x_sw),
    .io_x_sx(_2_28_io_x_sx),
    .io_x_sr(_2_28_io_x_sr),
    .io_x_pw(_2_28_io_x_pw),
    .io_x_px(_2_28_io_x_px),
    .io_x_pr(_2_28_io_x_pr),
    .io_x_pal(_2_28_io_x_pal),
    .io_x_paa(_2_28_io_x_paa),
    .io_x_eff(_2_28_io_x_eff),
    .io_x_c(_2_28_io_x_c),
    .io_y_ppn(_2_28_io_y_ppn),
    .io_y_u(_2_28_io_y_u),
    .io_y_ae(_2_28_io_y_ae),
    .io_y_sw(_2_28_io_y_sw),
    .io_y_sx(_2_28_io_y_sx),
    .io_y_sr(_2_28_io_y_sr),
    .io_y_pw(_2_28_io_y_pw),
    .io_y_px(_2_28_io_y_px),
    .io_y_pr(_2_28_io_y_pr),
    .io_y_pal(_2_28_io_y_pal),
    .io_y_paa(_2_28_io_y_paa),
    .io_y_eff(_2_28_io_y_eff),
    .io_y_c(_2_28_io_y_c)
  );
  _2_1 _2_29 (
    .io_x_ppn(_2_29_io_x_ppn),
    .io_x_u(_2_29_io_x_u),
    .io_x_ae(_2_29_io_x_ae),
    .io_x_sw(_2_29_io_x_sw),
    .io_x_sx(_2_29_io_x_sx),
    .io_x_sr(_2_29_io_x_sr),
    .io_x_pw(_2_29_io_x_pw),
    .io_x_px(_2_29_io_x_px),
    .io_x_pr(_2_29_io_x_pr),
    .io_x_pal(_2_29_io_x_pal),
    .io_x_paa(_2_29_io_x_paa),
    .io_x_eff(_2_29_io_x_eff),
    .io_x_c(_2_29_io_x_c),
    .io_y_ppn(_2_29_io_y_ppn),
    .io_y_u(_2_29_io_y_u),
    .io_y_ae(_2_29_io_y_ae),
    .io_y_sw(_2_29_io_y_sw),
    .io_y_sx(_2_29_io_y_sx),
    .io_y_sr(_2_29_io_y_sr),
    .io_y_pw(_2_29_io_y_pw),
    .io_y_px(_2_29_io_y_px),
    .io_y_pr(_2_29_io_y_pr),
    .io_y_pal(_2_29_io_y_pal),
    .io_y_paa(_2_29_io_y_paa),
    .io_y_eff(_2_29_io_y_eff),
    .io_y_c(_2_29_io_y_c)
  );
  _2_1 _2_30 (
    .io_x_ppn(_2_30_io_x_ppn),
    .io_x_u(_2_30_io_x_u),
    .io_x_ae(_2_30_io_x_ae),
    .io_x_sw(_2_30_io_x_sw),
    .io_x_sx(_2_30_io_x_sx),
    .io_x_sr(_2_30_io_x_sr),
    .io_x_pw(_2_30_io_x_pw),
    .io_x_px(_2_30_io_x_px),
    .io_x_pr(_2_30_io_x_pr),
    .io_x_pal(_2_30_io_x_pal),
    .io_x_paa(_2_30_io_x_paa),
    .io_x_eff(_2_30_io_x_eff),
    .io_x_c(_2_30_io_x_c),
    .io_y_ppn(_2_30_io_y_ppn),
    .io_y_u(_2_30_io_y_u),
    .io_y_ae(_2_30_io_y_ae),
    .io_y_sw(_2_30_io_y_sw),
    .io_y_sx(_2_30_io_y_sx),
    .io_y_sr(_2_30_io_y_sr),
    .io_y_pw(_2_30_io_y_pw),
    .io_y_px(_2_30_io_y_px),
    .io_y_pr(_2_30_io_y_pr),
    .io_y_pal(_2_30_io_y_pal),
    .io_y_paa(_2_30_io_y_paa),
    .io_y_eff(_2_30_io_y_eff),
    .io_y_c(_2_30_io_y_c)
  );
  _2_1 _2_31 (
    .io_x_ppn(_2_31_io_x_ppn),
    .io_x_u(_2_31_io_x_u),
    .io_x_ae(_2_31_io_x_ae),
    .io_x_sw(_2_31_io_x_sw),
    .io_x_sx(_2_31_io_x_sx),
    .io_x_sr(_2_31_io_x_sr),
    .io_x_pw(_2_31_io_x_pw),
    .io_x_px(_2_31_io_x_px),
    .io_x_pr(_2_31_io_x_pr),
    .io_x_pal(_2_31_io_x_pal),
    .io_x_paa(_2_31_io_x_paa),
    .io_x_eff(_2_31_io_x_eff),
    .io_x_c(_2_31_io_x_c),
    .io_y_ppn(_2_31_io_y_ppn),
    .io_y_u(_2_31_io_y_u),
    .io_y_ae(_2_31_io_y_ae),
    .io_y_sw(_2_31_io_y_sw),
    .io_y_sx(_2_31_io_y_sx),
    .io_y_sr(_2_31_io_y_sr),
    .io_y_pw(_2_31_io_y_pw),
    .io_y_px(_2_31_io_y_px),
    .io_y_pr(_2_31_io_y_pr),
    .io_y_pal(_2_31_io_y_pal),
    .io_y_paa(_2_31_io_y_paa),
    .io_y_eff(_2_31_io_y_eff),
    .io_y_c(_2_31_io_y_c)
  );
  _2_1 _2_32 (
    .io_x_ppn(_2_32_io_x_ppn),
    .io_x_u(_2_32_io_x_u),
    .io_x_ae(_2_32_io_x_ae),
    .io_x_sw(_2_32_io_x_sw),
    .io_x_sx(_2_32_io_x_sx),
    .io_x_sr(_2_32_io_x_sr),
    .io_x_pw(_2_32_io_x_pw),
    .io_x_px(_2_32_io_x_px),
    .io_x_pr(_2_32_io_x_pr),
    .io_x_pal(_2_32_io_x_pal),
    .io_x_paa(_2_32_io_x_paa),
    .io_x_eff(_2_32_io_x_eff),
    .io_x_c(_2_32_io_x_c),
    .io_y_ppn(_2_32_io_y_ppn),
    .io_y_u(_2_32_io_y_u),
    .io_y_ae(_2_32_io_y_ae),
    .io_y_sw(_2_32_io_y_sw),
    .io_y_sx(_2_32_io_y_sx),
    .io_y_sr(_2_32_io_y_sr),
    .io_y_pw(_2_32_io_y_pw),
    .io_y_px(_2_32_io_y_px),
    .io_y_pr(_2_32_io_y_pr),
    .io_y_pal(_2_32_io_y_pal),
    .io_y_paa(_2_32_io_y_paa),
    .io_y_eff(_2_32_io_y_eff),
    .io_y_c(_2_32_io_y_c)
  );
  _2_1 _2_33 (
    .io_x_ppn(_2_33_io_x_ppn),
    .io_x_u(_2_33_io_x_u),
    .io_x_ae(_2_33_io_x_ae),
    .io_x_sw(_2_33_io_x_sw),
    .io_x_sx(_2_33_io_x_sx),
    .io_x_sr(_2_33_io_x_sr),
    .io_x_pw(_2_33_io_x_pw),
    .io_x_px(_2_33_io_x_px),
    .io_x_pr(_2_33_io_x_pr),
    .io_x_pal(_2_33_io_x_pal),
    .io_x_paa(_2_33_io_x_paa),
    .io_x_eff(_2_33_io_x_eff),
    .io_x_c(_2_33_io_x_c),
    .io_y_ppn(_2_33_io_y_ppn),
    .io_y_u(_2_33_io_y_u),
    .io_y_ae(_2_33_io_y_ae),
    .io_y_sw(_2_33_io_y_sw),
    .io_y_sx(_2_33_io_y_sx),
    .io_y_sr(_2_33_io_y_sr),
    .io_y_pw(_2_33_io_y_pw),
    .io_y_px(_2_33_io_y_px),
    .io_y_pr(_2_33_io_y_pr),
    .io_y_pal(_2_33_io_y_pal),
    .io_y_paa(_2_33_io_y_paa),
    .io_y_eff(_2_33_io_y_eff),
    .io_y_c(_2_33_io_y_c)
  );
  _2_1 _2_34 (
    .io_x_ppn(_2_34_io_x_ppn),
    .io_x_u(_2_34_io_x_u),
    .io_x_ae(_2_34_io_x_ae),
    .io_x_sw(_2_34_io_x_sw),
    .io_x_sx(_2_34_io_x_sx),
    .io_x_sr(_2_34_io_x_sr),
    .io_x_pw(_2_34_io_x_pw),
    .io_x_px(_2_34_io_x_px),
    .io_x_pr(_2_34_io_x_pr),
    .io_x_pal(_2_34_io_x_pal),
    .io_x_paa(_2_34_io_x_paa),
    .io_x_eff(_2_34_io_x_eff),
    .io_x_c(_2_34_io_x_c),
    .io_y_ppn(_2_34_io_y_ppn),
    .io_y_u(_2_34_io_y_u),
    .io_y_ae(_2_34_io_y_ae),
    .io_y_sw(_2_34_io_y_sw),
    .io_y_sx(_2_34_io_y_sx),
    .io_y_sr(_2_34_io_y_sr),
    .io_y_pw(_2_34_io_y_pw),
    .io_y_px(_2_34_io_y_px),
    .io_y_pr(_2_34_io_y_pr),
    .io_y_pal(_2_34_io_y_pal),
    .io_y_paa(_2_34_io_y_paa),
    .io_y_eff(_2_34_io_y_eff),
    .io_y_c(_2_34_io_y_c)
  );
  _2_1 _2_35 (
    .io_x_ppn(_2_35_io_x_ppn),
    .io_x_u(_2_35_io_x_u),
    .io_x_ae(_2_35_io_x_ae),
    .io_x_sw(_2_35_io_x_sw),
    .io_x_sx(_2_35_io_x_sx),
    .io_x_sr(_2_35_io_x_sr),
    .io_x_pw(_2_35_io_x_pw),
    .io_x_px(_2_35_io_x_px),
    .io_x_pr(_2_35_io_x_pr),
    .io_x_pal(_2_35_io_x_pal),
    .io_x_paa(_2_35_io_x_paa),
    .io_x_eff(_2_35_io_x_eff),
    .io_x_c(_2_35_io_x_c),
    .io_y_ppn(_2_35_io_y_ppn),
    .io_y_u(_2_35_io_y_u),
    .io_y_ae(_2_35_io_y_ae),
    .io_y_sw(_2_35_io_y_sw),
    .io_y_sx(_2_35_io_y_sx),
    .io_y_sr(_2_35_io_y_sr),
    .io_y_pw(_2_35_io_y_pw),
    .io_y_px(_2_35_io_y_px),
    .io_y_pr(_2_35_io_y_pr),
    .io_y_pal(_2_35_io_y_pal),
    .io_y_paa(_2_35_io_y_paa),
    .io_y_eff(_2_35_io_y_eff),
    .io_y_c(_2_35_io_y_c)
  );
  _2_1 _2_36 (
    .io_x_ppn(_2_36_io_x_ppn),
    .io_x_u(_2_36_io_x_u),
    .io_x_ae(_2_36_io_x_ae),
    .io_x_sw(_2_36_io_x_sw),
    .io_x_sx(_2_36_io_x_sx),
    .io_x_sr(_2_36_io_x_sr),
    .io_x_pw(_2_36_io_x_pw),
    .io_x_px(_2_36_io_x_px),
    .io_x_pr(_2_36_io_x_pr),
    .io_x_pal(_2_36_io_x_pal),
    .io_x_paa(_2_36_io_x_paa),
    .io_x_eff(_2_36_io_x_eff),
    .io_x_c(_2_36_io_x_c),
    .io_y_ppn(_2_36_io_y_ppn),
    .io_y_u(_2_36_io_y_u),
    .io_y_ae(_2_36_io_y_ae),
    .io_y_sw(_2_36_io_y_sw),
    .io_y_sx(_2_36_io_y_sx),
    .io_y_sr(_2_36_io_y_sr),
    .io_y_pw(_2_36_io_y_pw),
    .io_y_px(_2_36_io_y_px),
    .io_y_pr(_2_36_io_y_pr),
    .io_y_pal(_2_36_io_y_pal),
    .io_y_paa(_2_36_io_y_paa),
    .io_y_eff(_2_36_io_y_eff),
    .io_y_c(_2_36_io_y_c)
  );
  _2_1 _2_37 (
    .io_x_ppn(_2_37_io_x_ppn),
    .io_x_u(_2_37_io_x_u),
    .io_x_ae(_2_37_io_x_ae),
    .io_x_sw(_2_37_io_x_sw),
    .io_x_sx(_2_37_io_x_sx),
    .io_x_sr(_2_37_io_x_sr),
    .io_x_pw(_2_37_io_x_pw),
    .io_x_px(_2_37_io_x_px),
    .io_x_pr(_2_37_io_x_pr),
    .io_x_pal(_2_37_io_x_pal),
    .io_x_paa(_2_37_io_x_paa),
    .io_x_eff(_2_37_io_x_eff),
    .io_x_c(_2_37_io_x_c),
    .io_y_ppn(_2_37_io_y_ppn),
    .io_y_u(_2_37_io_y_u),
    .io_y_ae(_2_37_io_y_ae),
    .io_y_sw(_2_37_io_y_sw),
    .io_y_sx(_2_37_io_y_sx),
    .io_y_sr(_2_37_io_y_sr),
    .io_y_pw(_2_37_io_y_pw),
    .io_y_px(_2_37_io_y_px),
    .io_y_pr(_2_37_io_y_pr),
    .io_y_pal(_2_37_io_y_pal),
    .io_y_paa(_2_37_io_y_paa),
    .io_y_eff(_2_37_io_y_eff),
    .io_y_c(_2_37_io_y_c)
  );
  _2_1 _2_38 (
    .io_x_ppn(_2_38_io_x_ppn),
    .io_x_u(_2_38_io_x_u),
    .io_x_ae(_2_38_io_x_ae),
    .io_x_sw(_2_38_io_x_sw),
    .io_x_sx(_2_38_io_x_sx),
    .io_x_sr(_2_38_io_x_sr),
    .io_x_pw(_2_38_io_x_pw),
    .io_x_px(_2_38_io_x_px),
    .io_x_pr(_2_38_io_x_pr),
    .io_x_pal(_2_38_io_x_pal),
    .io_x_paa(_2_38_io_x_paa),
    .io_x_eff(_2_38_io_x_eff),
    .io_x_c(_2_38_io_x_c),
    .io_y_ppn(_2_38_io_y_ppn),
    .io_y_u(_2_38_io_y_u),
    .io_y_ae(_2_38_io_y_ae),
    .io_y_sw(_2_38_io_y_sw),
    .io_y_sx(_2_38_io_y_sx),
    .io_y_sr(_2_38_io_y_sr),
    .io_y_pw(_2_38_io_y_pw),
    .io_y_px(_2_38_io_y_px),
    .io_y_pr(_2_38_io_y_pr),
    .io_y_pal(_2_38_io_y_pal),
    .io_y_paa(_2_38_io_y_paa),
    .io_y_eff(_2_38_io_y_eff),
    .io_y_c(_2_38_io_y_c)
  );

`define MY_ASSIGNMENT
`ifdef MY_ASSIGNMENT
  assign priv_s = io_ptw_status_dprv[0];
  assign priv_uses_vm = io_ptw_status_dprv <= 2'h1; 

  assign vm_enabled = io_ptw_ptbr_mode & priv_uses_vm & !io_req_bits_passthrough;

  assign vpn = io_req_bits_vaddr[31:12];

  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0];

  wire _T_4 = state == 2'h1;
  assign invalidate_refill = _T_4 | (state == 2'h3);

  wire _T_25 = special_entry_level < 1'h1;
  wire [19:0] _T_27 = _T_25 ? vpn : 20'h0;
  assign mpu_ppn = io_ptw_resp_valid ? refill_ppn 
		: vm_enabled ? {_2_io_y_ppn[19:10], (_T_27[9:0] | _2_io_y_ppn[9:0])} 
		: io_req_bits_vaddr[31:12];

  assign mpu_physaddr = {mpu_ppn, io_req_bits_vaddr[11:0]};

  assign mpu_priv = (io_ptw_resp_valid | io_req_bits_passthrough) ? 3'h1 : {io_ptw_status_debug,io_ptw_status_dprv};

  wire [32:0] _T_48 = {1'b0,$signed(mpu_physaddr ^ 32'h2000000)};
  wire [32:0] _T_53 = {1'b0,$signed(mpu_physaddr)};
  wire _T_56 = $signed($signed(_T_53) & $signed(-33'sh1000)) == $signed(33'sh0);
  wire [32:0] _T_63 = {1'b0,$signed(mpu_physaddr ^ 32'h80000000)};
  assign legal_address = ($signed($signed({1'b0,$signed(mpu_physaddr ^ 32'h3000)}) & $signed(-33'sh1000)) == $signed(33'sh0)) 
			| ($signed($signed({1'b0,$signed(mpu_physaddr ^ 32'hc000000)}) & $signed(-33'sh4000000)) == $signed(33'sh0)) 
			| ($signed($signed(_T_48) & $signed(-33'sh10000)) == $signed(33'sh0)) 
			| _T_56 
			| ($signed($signed({1'b0,$signed(mpu_physaddr ^ 32'h10000)}) & $signed(-33'sh10000)) == $signed(33'sh0)) 
			| ($signed($signed(_T_63) & $signed(-33'sh10000000)) == $signed(33'sh0)) 
			| ($signed($signed({1'b0,$signed(mpu_physaddr ^ 32'h60000000)}) & $signed(-33'sh20000000)) == $signed(33'sh0));

  assign cacheable = legal_address & ($signed($signed(_T_63) & $signed(33'sh80000000)) == $signed(33'sh0));

  assign deny_access_to_debug = (mpu_priv <= 3'h3) & ($signed($signed(_T_53) & $signed(-33'sh1000)) == $signed(33'sh0));

  wire _T_197 = deny_access_to_debug == 1'h0;
  assign prot_r = legal_address & _T_197 & pmp_io_r;

  wire _T_146 = $signed($signed({1'b0,$signed(mpu_physaddr ^ 32'h8000000)}) & $signed(33'shc8000000)) == $signed(33'sh0);
  wire _T_172 = ($signed($signed(_T_53) & $signed(33'shc8010000)) == $signed(33'sh0)) 
		| _T_146;
  wire _T_213 = $signed($signed({1'b0,$signed(mpu_physaddr ^ 32'h80000000)}) & $signed(33'shc0000000)) == $signed(33'sh0);
  wire _T_218 = $signed($signed({1'b0,$signed(mpu_physaddr ^ 32'h40000000)}) & $signed(33'shc0000000)) == $signed(33'sh0);
  assign prot_w = (legal_address & 
			( _T_172 
			| _T_213 
			| _T_218)
			 & _T_197) & pmp_io_w;
// Passed
  assign prot_al = legal_address & _T_172;

  assign prot_x = legal_address & 
			(($signed($signed(_T_53) & $signed(33'shca000000)) == $signed(33'sh0)) 
			| _T_213 
			| _T_218) 
			& _T_197 & pmp_io_x;

  assign prot_eff = legal_address & 
			(_T_146 
			| ($signed($signed({1'b0,$signed(mpu_physaddr ^ 32'h2000000)}) & $signed(33'shca010000)) == $signed(33'sh0)) 
			| ($signed($signed(_T_53) & $signed(33'shca012000)) == $signed(33'sh0)) 
			| _T_218);

  wire _T_379 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1 | sectored_entries_0_valid_2 | sectored_entries_0_valid_3;
  wire [19:0] _T_380 = sectored_entries_0_tag ^ vpn;
  wire _T_382 = _T_380[19:2] == 18'h0;
  assign sector_hits_0 = _T_379 & _T_382;

  wire _T_385 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1 | sectored_entries_1_valid_2 | sectored_entries_1_valid_3;
  wire [19:0] _T_386 = sectored_entries_1_tag ^ vpn;
  wire _T_388 = _T_386[19:2] == 18'h0; 
  assign sector_hits_1 = _T_385 & _T_388;

  wire _T_391 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1 | sectored_entries_2_valid_2 | sectored_entries_2_valid_3;
  wire [19:0] _T_392 = sectored_entries_2_tag ^ vpn;
  wire _T_394 = _T_392[19:2] == 18'h0;
  assign sector_hits_2 = _T_391 & _T_394;

  wire _T_397 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1 | sectored_entries_3_valid_2 | sectored_entries_3_valid_3;
  wire [19:0] _T_398 = sectored_entries_3_tag ^ vpn;
  wire _T_400 = _T_398[19:2] == 18'h0;
  assign sector_hits_3 = _T_397 & _T_400;

  wire _T_403 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1 | sectored_entries_4_valid_2 | sectored_entries_4_valid_3;
  wire [19:0] _T_404 = sectored_entries_4_tag ^ vpn;
  wire _T_406 = _T_404[19:2] == 18'h0;
  assign sector_hits_4 = _T_403 & _T_406;

  wire _T_409 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1 | sectored_entries_5_valid_2 | sectored_entries_5_valid_3;
  wire [19:0] _T_410 = sectored_entries_5_tag ^ vpn;
  wire _T_412 = _T_410[19:2] == 18'h0;
  assign sector_hits_5 = _T_409 & _T_412;

  wire _T_415 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1 | sectored_entries_6_valid_2 | sectored_entries_6_valid_3;
  wire [19:0] _T_416 = sectored_entries_6_tag ^ vpn;
  wire _T_418 = _T_416[19:2] == 18'h0;
  assign sector_hits_6 = _T_415 & _T_418;

  wire _T_421 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1 | sectored_entries_7_valid_2 | sectored_entries_7_valid_3;
  wire [19:0] _T_422 = sectored_entries_7_tag ^ vpn;
  wire _T_424 = _T_422[19:2] == 18'h0;
  assign sector_hits_7 = _T_421 & _T_424;
// Passed
  assign superpage_hits_0 = superpage_entries_0_valid_0 & (superpage_entries_0_tag[19:10] == vpn[19:10]);

  assign superpage_hits_1 = superpage_entries_1_valid_0 & (superpage_entries_1_tag[19:10] == vpn[19:10]);

  assign superpage_hits_2 = superpage_entries_2_valid_0 & (superpage_entries_2_tag[19:10] == vpn[19:10]);

  assign superpage_hits_3 = superpage_entries_3_valid_0 & (superpage_entries_3_tag[19:10] == vpn[19:10]);

  wire [1:0] _T_477 = vpn[1:0];
  assign hitsVec_0 = vm_enabled & (2'h3 == _T_477 ? sectored_entries_0_valid_3 
				: 2'h2 == _T_477 ? sectored_entries_0_valid_2 
				: 2'h1 == _T_477 ? sectored_entries_0_valid_1 
				: sectored_entries_0_valid_0) & _T_382;

  assign hitsVec_1 = vm_enabled & (2'h3 == _T_477 ? sectored_entries_1_valid_3 
				: 2'h2 == _T_477 ? sectored_entries_1_valid_2 
				: 2'h1 == _T_477 ? sectored_entries_1_valid_1 
				: sectored_entries_1_valid_0) & _T_388;

  assign hitsVec_2 = vm_enabled & (2'h3 == _T_477 ? sectored_entries_2_valid_3 
				: 2'h2 == _T_477 ? sectored_entries_2_valid_2 
				: 2'h1 == _T_477 ? sectored_entries_2_valid_1 
				: sectored_entries_2_valid_0) & _T_394;

  assign hitsVec_3 = vm_enabled & (2'h3 == _T_477 ? sectored_entries_3_valid_3 
				: 2'h2 == _T_477 ? sectored_entries_3_valid_2 
				: 2'h1 == _T_477 ? sectored_entries_3_valid_1 
				: sectored_entries_3_valid_0) & _T_400;

  assign hitsVec_4 = vm_enabled & (2'h3 == _T_477 ? sectored_entries_4_valid_3 
				: 2'h2 == _T_477 ? sectored_entries_4_valid_2 
				: 2'h1 == _T_477 ? sectored_entries_4_valid_1 
				: sectored_entries_4_valid_0) & _T_406;

  assign hitsVec_5 = vm_enabled & (2'h3 == _T_477 ? sectored_entries_5_valid_3 
				: 2'h2 == _T_477 ? sectored_entries_5_valid_2 
				: 2'h1 == _T_477 ? sectored_entries_5_valid_1 
				: sectored_entries_5_valid_0) & _T_412;

  assign hitsVec_6 = vm_enabled & (2'h3 == _T_477 ? sectored_entries_6_valid_3 
				: 2'h2 == _T_477 ? sectored_entries_6_valid_2 
				: 2'h1 == _T_477 ? sectored_entries_6_valid_1 
				: sectored_entries_6_valid_0) & _T_418;

  assign hitsVec_7 = vm_enabled & (2'h3 == _T_477 ? sectored_entries_7_valid_3 
				: 2'h2 == _T_477 ? sectored_entries_7_valid_2 
				: 2'h1 == _T_477 ? sectored_entries_7_valid_1 
				: sectored_entries_7_valid_0) & _T_424;

  assign hitsVec_8 = vm_enabled & superpage_hits_0;
  assign hitsVec_9 = vm_enabled & superpage_hits_1;
  assign hitsVec_10 = vm_enabled & superpage_hits_2;
  assign hitsVec_11 = vm_enabled & superpage_hits_3;

  wire _T_586 = special_entry_valid_0 & (special_entry_tag[19:10] == vpn[19:10]) & ((special_entry_level < 1'h1) | (special_entry_tag[9:0] == vpn[9:0]));
  assign hitsVec_12 = vm_enabled & _T_586;

  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0};

  wire _T_598 = vm_enabled == 1'h0;
  assign hits = {_T_598,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0};

  assign ppn = (hitsVec_0 ? _2_1_io_y_ppn : 20'h0) 
  		| (hitsVec_1 ? _2_2_io_y_ppn : 20'h0)
  		| (hitsVec_2 ? _2_3_io_y_ppn : 20'h0)
  		| (hitsVec_3 ? _2_4_io_y_ppn : 20'h0)
  		| (hitsVec_4 ? _2_5_io_y_ppn : 20'h0)
  		| (hitsVec_5 ? _2_6_io_y_ppn : 20'h0)
  		| (hitsVec_6 ? _2_7_io_y_ppn : 20'h0)
  		| (hitsVec_7 ? _2_8_io_y_ppn : 20'h0)
  		| (hitsVec_8 ? {_2_9_io_y_ppn[19:10], (vpn[9:0] | _2_9_io_y_ppn[9:0])} : 20'h0)
  		| (hitsVec_9 ? {_2_10_io_y_ppn[19:10], (vpn[9:0] | _2_10_io_y_ppn[9:0])} : 20'h0)
  		| (hitsVec_10 ? {_2_11_io_y_ppn[19:10], (vpn[9:0] | _2_11_io_y_ppn[9:0])} : 20'h0)
  		| (hitsVec_11 ? {_2_12_io_y_ppn[19:10], (vpn[9:0] | _2_12_io_y_ppn[9:0])} : 20'h0)
  		| (hitsVec_12 ? {_2_13_io_y_ppn[19:10], (_T_27[9:0] | _2_13_io_y_ppn[9:0])} : 20'h0)
  		| (_T_598 ? vpn : 20'h0);

  assign ptw_ae_array = {1'h0,_2_26_io_y_ae,_2_25_io_y_ae,_2_24_io_y_ae,_2_23_io_y_ae,_2_22_io_y_ae,_2_21_io_y_ae,_2_20_io_y_ae,_2_19_io_y_ae,_2_18_io_y_ae,_2_17_io_y_ae,_2_16_io_y_ae,_2_15_io_y_ae,_2_14_io_y_ae};

  assign priv_rw_ok = ((!priv_s | io_ptw_status_sum) ? {_2_26_io_y_u,_2_25_io_y_u,_2_24_io_y_u,_2_23_io_y_u,_2_22_io_y_u,_2_21_io_y_u,_2_20_io_y_u,_2_19_io_y_u,_2_18_io_y_u,_2_17_io_y_u,_2_16_io_y_u,_2_15_io_y_u,_2_14_io_y_u} : 13'h0) 
			| (priv_s ? ~ {_2_26_io_y_u,_2_25_io_y_u,_2_24_io_y_u,_2_23_io_y_u,_2_22_io_y_u,_2_21_io_y_u,_2_20_io_y_u,_2_19_io_y_u,_2_18_io_y_u,_2_17_io_y_u,_2_16_io_y_u,_2_15_io_y_u,_2_14_io_y_u} : 13'h0);

  wire [12:0] _T_1663 = priv_rw_ok & ({_2_26_io_y_sr,_2_25_io_y_sr,_2_24_io_y_sr,_2_23_io_y_sr,_2_22_io_y_sr,_2_21_io_y_sr,_2_20_io_y_sr,_2_19_io_y_sr,_2_18_io_y_sr,_2_17_io_y_sr,_2_16_io_y_sr,_2_15_io_y_sr,_2_14_io_y_sr} | (io_ptw_status_mxr ? {_2_26_io_y_sx,_2_25_io_y_sx,_2_24_io_y_sx,_2_23_io_y_sx,_2_22_io_y_sx,_2_21_io_y_sx,_2_20_io_y_sx,_2_19_io_y_sx,_2_18_io_y_sx,_2_17_io_y_sx,_2_16_io_y_sx,_2_15_io_y_sx,_2_14_io_y_sx} : 13'h0));
  assign r_array = {1'h1,_T_1663};
// Passed
  wire [12:0] _T_1676 = priv_rw_ok & {_2_26_io_y_sw,_2_25_io_y_sw,_2_24_io_y_sw,_2_23_io_y_sw,_2_22_io_y_sw,_2_21_io_y_sw,_2_20_io_y_sw,_2_19_io_y_sw,_2_18_io_y_sw,_2_17_io_y_sw,_2_16_io_y_sw,_2_15_io_y_sw,_2_14_io_y_sw};
  assign w_array = {1'h1,_T_1676};

  wire [1:0] _T_1691 = prot_r ? 2'h3 : 2'h0;
  assign pr_array = {_T_1691,_2_38_io_y_pr,_2_37_io_y_pr,_2_36_io_y_pr,_2_35_io_y_pr,_2_34_io_y_pr,_2_33_io_y_pr,_2_32_io_y_pr,_2_31_io_y_pr,_2_30_io_y_pr,_2_29_io_y_pr,_2_28_io_y_pr,_2_27_io_y_pr} & (~ ptw_ae_array);

  wire [1:0] _T_1706 = prot_w ? 2'h3 : 2'h0;
  assign pw_array = {_T_1706,_2_38_io_y_pw,_2_37_io_y_pw,_2_36_io_y_pw,_2_35_io_y_pw,_2_34_io_y_pw,_2_33_io_y_pw,_2_32_io_y_pw,_2_31_io_y_pw,_2_30_io_y_pw,_2_29_io_y_pw,_2_28_io_y_pw,_2_27_io_y_pw} & (~ ptw_ae_array);

  wire [1:0] _T_1736 = prot_eff ? 2'h3 : 2'h0;
  assign eff_array = {_T_1736,_2_38_io_y_eff,_2_37_io_y_eff,_2_36_io_y_eff,_2_35_io_y_eff,_2_34_io_y_eff,_2_33_io_y_eff,_2_32_io_y_eff,_2_31_io_y_eff,_2_30_io_y_eff,_2_29_io_y_eff,_2_28_io_y_eff,_2_27_io_y_eff};

  wire [1:0] _T_1749 = cacheable ? 2'h3 : 2'h0;
  assign c_array = {_T_1749,_2_38_io_y_c,_2_37_io_y_c,_2_36_io_y_c,_2_35_io_y_c,_2_34_io_y_c,_2_33_io_y_c,_2_32_io_y_c,_2_31_io_y_c,_2_30_io_y_c,_2_29_io_y_c,_2_28_io_y_c,_2_27_io_y_c};

  wire [1:0] _T_1762 = prot_al ? 2'h3 : 2'h0;
  assign paa_array = {_T_1762,_2_38_io_y_paa,_2_37_io_y_paa,_2_36_io_y_paa,_2_35_io_y_paa,_2_34_io_y_paa,_2_33_io_y_paa,_2_32_io_y_paa,_2_31_io_y_paa,_2_30_io_y_paa,_2_29_io_y_paa,_2_28_io_y_paa,_2_27_io_y_paa};

  assign pal_array = {_T_1762,_2_38_io_y_pal,_2_37_io_y_pal,_2_36_io_y_pal,_2_35_io_y_pal,_2_34_io_y_pal,_2_33_io_y_pal,_2_32_io_y_pal,_2_31_io_y_pal,_2_30_io_y_pal,_2_29_io_y_pal,_2_28_io_y_pal,_2_27_io_y_pal};

  assign paa_array_if_cached = paa_array | c_array;
  assign pal_array_if_cached = pal_array | c_array;

  wire [3:0] _T_1804 = (4'h1 << io_req_bits_size) - 4'h1;
  assign misaligned = (io_req_bits_vaddr & {{28'd0}, _T_1804}) != 32'h0;

  wire _T_1806 = io_req_bits_cmd == 5'h6;
  wire _T_1807 = io_req_bits_cmd == 5'h7;
  assign cmd_lrsc = _T_1806 | _T_1807;

  assign cmd_amo_logical = (io_req_bits_cmd == 5'h4) 
				| (io_req_bits_cmd == 5'h9) 
				| (io_req_bits_cmd == 5'ha) 
				| (io_req_bits_cmd == 5'hb);

  assign cmd_amo_arithmetic = (io_req_bits_cmd == 5'h8) 
				| (io_req_bits_cmd == 5'hc) 
				| (io_req_bits_cmd == 5'hd) 
				| (io_req_bits_cmd == 5'he) 
				| (io_req_bits_cmd == 5'hf);
// Passed
  wire _T_1846 = cmd_amo_logical | cmd_amo_arithmetic;
  assign cmd_read = (io_req_bits_cmd == 5'h0) 
			| (io_req_bits_cmd == 5'h6) 
			| _T_1807 
			| _T_1846;

  assign cmd_write = (io_req_bits_cmd == 5'h1) 
			| (io_req_bits_cmd == 5'h11) 
			| _T_1807 
			| _T_1846;

  assign cmd_write_perms = cmd_write 
			| (io_req_bits_cmd == 5'h5) 
			| (io_req_bits_cmd == 5'h17);

  assign ae_array = (misaligned ? eff_array : 14'h0) 
			| (cmd_lrsc ? (~ c_array) : 14'h0);

  assign ae_ld_array = cmd_read ? (ae_array | (~ pr_array)) : 14'h0;

  assign ae_st_array = (cmd_write_perms ? (ae_array | (~ pw_array)) : 14'h0) 
			| (cmd_amo_logical ? ~ pal_array_if_cached : 14'h0) 
			| (cmd_amo_arithmetic ? ~ paa_array_if_cached : 14'h0);

  assign ma_ld_array = (misaligned & cmd_read) ? (~ eff_array) : 14'h0;

  assign ma_st_array = (misaligned & cmd_write) ? (~ eff_array) : 14'h0;

  assign pf_ld_array = cmd_read ? (~ (r_array | ptw_ae_array)) : 14'h0;

  assign pf_st_array = cmd_write_perms ? (~ (w_array | ptw_ae_array)) : 14'h0;

  assign tlb_hit = real_hits != 13'h0;

  assign tlb_miss = vm_enabled & !tlb_hit;

  wire _T_1995 = real_hits[0];
  wire _T_1998 = real_hits[1];
  wire _T_2000 = real_hits[2];
  wire _T_2011 = real_hits[3];
  wire _T_2014 = real_hits[4];
  wire _T_2016 = real_hits[5];
  wire _T_2032 = real_hits[6];
  wire _T_2035 = real_hits[7];
  wire _T_2037 = real_hits[8];
  wire _T_2049 = real_hits[9];
  wire _T_2051 = real_hits[10];
  wire _T_2058 = real_hits[11];
  wire _T_2060 = real_hits[12];
  assign multipleHits = (real_hits[1] & real_hits[2]) 
			| (real_hits[0] & (real_hits[1] | real_hits[2])) 
			| (real_hits[4] & real_hits[5]) 
			| (real_hits[0] & (real_hits[4] | real_hits[5]))
			| ((_T_1995 | _T_1998 | _T_2000) & (_T_2011 | _T_2014 | _T_2016)) 
			| (_T_2035 & _T_2037) 
			| (_T_2032 & (_T_2035 | _T_2037)) 
			| (_T_2049 & _T_2051) 
			| (_T_2058 & _T_2060) 
			| ((_T_2049 | _T_2051) & (_T_2058 | _T_2060)) 
			| ((_T_2032 | _T_2035 | _T_2037) & (_T_2049 | _T_2051 | _T_2058 | _T_2060)) 
			| ((_T_1995 | _T_1998 | _T_2000 | _T_2011 | _T_2014 | _T_2016) & (_T_2032 | _T_2035 | _T_2037 | _T_2049 | _T_2051 | _T_2058 | _T_2060));
// Passed
  assign io_req_ready = state == 2'h0;

  assign io_resp_miss = io_ptw_resp_valid | tlb_miss | multipleHits;

  assign io_resp_paddr = {ppn, io_req_bits_vaddr[11:0]};

  assign io_resp_pf_ld = (pf_ld_array & hits) != 14'h0;

  assign io_resp_pf_st = (pf_st_array & hits) != 14'h0;

  assign io_resp_ae_ld = (ae_ld_array & hits) != 14'h0;

  assign io_resp_ae_st = (ae_st_array & hits) != 14'h0;
  assign io_resp_ma_ld = (ma_ld_array & hits) != 14'h0;
  assign io_resp_ma_st = (ma_st_array & hits) != 14'h0;
  assign io_resp_cacheable = (c_array & hits) != 14'h0;
  assign io_ptw_req_valid = state == 2'h1;
  assign io_ptw_req_bits_bits_addr = r_refill_tag;

  assign _2_io_x_ppn = special_entry_data_0[33:14];
  assign _2_io_x_u = special_entry_data_0[13];
  assign _2_io_x_ae = special_entry_data_0[11];
  assign _2_io_x_sw = special_entry_data_0[10];
  assign _2_io_x_sx = special_entry_data_0[9]; 
  assign _2_io_x_sr = special_entry_data_0[8]; 
  assign _2_io_x_pw = special_entry_data_0[7]; 
  assign _2_io_x_px = special_entry_data_0[6]; 
  assign _2_io_x_pr = special_entry_data_0[5]; 
  assign _2_io_x_pal = special_entry_data_0[4];
  assign _2_io_x_paa = special_entry_data_0[3];
  assign _2_io_x_eff = special_entry_data_0[2];
  assign _2_io_x_c = special_entry_data_0[1]; 

  assign pmp_io_prv = mpu_priv[1:0];
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr;
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask;
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr;
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask;
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr;
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask;
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr;
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask;
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr;
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask;
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr;
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask;
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr;
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask;
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr;
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask;
  assign pmp_io_addr = {mpu_ppn, io_req_bits_vaddr[11:0]};

  wire [33:0] _GEN_35 = 2'h3 == _T_477 ? sectored_entries_0_data_3 
		: 2'h2 == _T_477 ? sectored_entries_0_data_2 
		: 2'h1 == _T_477 ? sectored_entries_0_data_1 
		: sectored_entries_0_data_0;
  assign _2_1_io_x_ppn = _GEN_35[33:14];
  assign _2_1_io_x_u = _GEN_35[13];
  assign _2_1_io_x_ae = _GEN_35[11];
  assign _2_1_io_x_sw = _GEN_35[10];
  assign _2_1_io_x_sx = _GEN_35[9];
  assign _2_1_io_x_sr = _GEN_35[8];
  assign _2_1_io_x_pw = _GEN_35[7];
  assign _2_1_io_x_px = _GEN_35[6];
  assign _2_1_io_x_pr = _GEN_35[5];
  assign _2_1_io_x_pal = _GEN_35[4];
  assign _2_1_io_x_paa = _GEN_35[3];
  assign _2_1_io_x_eff = _GEN_35[2];
  assign _2_1_io_x_c = _GEN_35[1];

  wire [33:0] _GEN_39 = 2'h3 == _T_477 ? sectored_entries_1_data_3 
		: 2'h2 == _T_477 ? sectored_entries_1_data_2 
		: 2'h1 == _T_477 ? sectored_entries_1_data_1 
		: sectored_entries_1_data_0;
  assign _2_2_io_x_ppn = _GEN_39[33:14];
  assign _2_2_io_x_u = _GEN_39[13];
  assign _2_2_io_x_ae = _GEN_39[11];
  assign _2_2_io_x_sw = _GEN_39[10];
  assign _2_2_io_x_sx = _GEN_39[9];
  assign _2_2_io_x_sr = _GEN_39[8];
  assign _2_2_io_x_pw = _GEN_39[7];
  assign _2_2_io_x_px = _GEN_39[6];
  assign _2_2_io_x_pr = _GEN_39[5];
  assign _2_2_io_x_pal = _GEN_39[4];
  assign _2_2_io_x_paa = _GEN_39[3];
  assign _2_2_io_x_eff = _GEN_39[2];
  assign _2_2_io_x_c = _GEN_39[1];

  wire [33:0] _GEN_43 = 2'h3 == _T_477 ? sectored_entries_2_data_3 
		: 2'h2 == _T_477 ? sectored_entries_2_data_2 
		: 2'h1 == _T_477 ? sectored_entries_2_data_1 
		: sectored_entries_2_data_0;
  assign _2_3_io_x_ppn = _GEN_43[33:14];
  assign _2_3_io_x_u = _GEN_43[13];
  assign _2_3_io_x_ae = _GEN_43[11];
  assign _2_3_io_x_sw = _GEN_43[10];
  assign _2_3_io_x_sx = _GEN_43[9]; 
  assign _2_3_io_x_sr = _GEN_43[8]; 
  assign _2_3_io_x_pw = _GEN_43[7]; 
  assign _2_3_io_x_px = _GEN_43[6]; 
  assign _2_3_io_x_pr = _GEN_43[5]; 
  assign _2_3_io_x_pal = _GEN_43[4];
  assign _2_3_io_x_paa = _GEN_43[3];
  assign _2_3_io_x_eff = _GEN_43[2];
  assign _2_3_io_x_c = _GEN_43[1];

  wire [33:0] _GEN_47 = 2'h3 == _T_477 ? sectored_entries_3_data_3 
		: 2'h2 == _T_477 ? sectored_entries_3_data_2 
		: 2'h1 == _T_477 ? sectored_entries_3_data_1 
		: sectored_entries_3_data_0;
  assign _2_4_io_x_ppn = _GEN_47[33:14];
  assign _2_4_io_x_u = _GEN_47[13]; 
  assign _2_4_io_x_ae = _GEN_47[11];
  assign _2_4_io_x_sw = _GEN_47[10];
  assign _2_4_io_x_sx = _GEN_47[9]; 
  assign _2_4_io_x_sr = _GEN_47[8]; 
  assign _2_4_io_x_pw = _GEN_47[7]; 
  assign _2_4_io_x_px = _GEN_47[6]; 
  assign _2_4_io_x_pr = _GEN_47[5]; 
  assign _2_4_io_x_pal = _GEN_47[4];
  assign _2_4_io_x_paa = _GEN_47[3];
  assign _2_4_io_x_eff = _GEN_47[2];
  assign _2_4_io_x_c = _GEN_47[1]; 

  wire [33:0] _GEN_51 = 2'h3 == _T_477 ? sectored_entries_4_data_3 
		: 2'h2 == _T_477 ? sectored_entries_4_data_2 
		: 2'h1 == _T_477 ? sectored_entries_4_data_1 
		: sectored_entries_4_data_0; 
  assign _2_5_io_x_ppn = _GEN_51[33:14];
  assign _2_5_io_x_u = _GEN_51[13]; 
  assign _2_5_io_x_ae = _GEN_51[11];
  assign _2_5_io_x_sw = _GEN_51[10];
  assign _2_5_io_x_sx = _GEN_51[9]; 
  assign _2_5_io_x_sr = _GEN_51[8]; 
  assign _2_5_io_x_pw = _GEN_51[7]; 
  assign _2_5_io_x_px = _GEN_51[6]; 
  assign _2_5_io_x_pr = _GEN_51[5]; 
  assign _2_5_io_x_pal = _GEN_51[4];
  assign _2_5_io_x_paa = _GEN_51[3];
  assign _2_5_io_x_eff = _GEN_51[2];
  assign _2_5_io_x_c = _GEN_51[1]; 

  wire [33:0] _GEN_55 = 2'h3 == _T_477 ? sectored_entries_5_data_3 
		: 2'h2 == _T_477 ? sectored_entries_5_data_2 
		: 2'h1 == _T_477 ? sectored_entries_5_data_1 
		: sectored_entries_5_data_0;
  assign _2_6_io_x_ppn = _GEN_55[33:14];
  assign _2_6_io_x_u = _GEN_55[13]; 
  assign _2_6_io_x_ae = _GEN_55[11];
  assign _2_6_io_x_sw = _GEN_55[10];
  assign _2_6_io_x_sx = _GEN_55[9]; 
  assign _2_6_io_x_sr = _GEN_55[8]; 
  assign _2_6_io_x_pw = _GEN_55[7]; 
  assign _2_6_io_x_px = _GEN_55[6]; 
  assign _2_6_io_x_pr = _GEN_55[5]; 
  assign _2_6_io_x_pal = _GEN_55[4];
  assign _2_6_io_x_paa = _GEN_55[3];
  assign _2_6_io_x_eff = _GEN_55[2];
  assign _2_6_io_x_c = _GEN_55[1]; 

  wire [33:0] _GEN_59 = 2'h3 == _T_477 ? sectored_entries_6_data_3 
		: 2'h2 == _T_477 ? sectored_entries_6_data_2 
		: 2'h1 == _T_477 ? sectored_entries_6_data_1 
		: sectored_entries_6_data_0;
  assign _2_7_io_x_ppn = _GEN_59[33:14];
  assign _2_7_io_x_u = _GEN_59[13]; 
  assign _2_7_io_x_ae = _GEN_59[11];
  assign _2_7_io_x_sw = _GEN_59[10];
  assign _2_7_io_x_sx = _GEN_59[9]; 
  assign _2_7_io_x_sr = _GEN_59[8]; 
  assign _2_7_io_x_pw = _GEN_59[7]; 
  assign _2_7_io_x_px = _GEN_59[6]; 
  assign _2_7_io_x_pr = _GEN_59[5]; 
  assign _2_7_io_x_pal = _GEN_59[4];
  assign _2_7_io_x_paa = _GEN_59[3];
  assign _2_7_io_x_eff = _GEN_59[2];
  assign _2_7_io_x_c = _GEN_59[1]; 

  wire [33:0] _GEN_63 = 2'h3 == _T_477 ? sectored_entries_7_data_3 
		: 2'h2 == _T_477 ? sectored_entries_7_data_2 
		: 2'h1 == _T_477 ? sectored_entries_7_data_1 
		: sectored_entries_7_data_0;
  assign _2_8_io_x_ppn = _GEN_63[33:14];
  assign _2_8_io_x_u = _GEN_63[13]; 
  assign _2_8_io_x_ae = _GEN_63[11];
  assign _2_8_io_x_sw = _GEN_63[10];
  assign _2_8_io_x_sx = _GEN_63[9]; 
  assign _2_8_io_x_sr = _GEN_63[8]; 
  assign _2_8_io_x_pw = _GEN_63[7]; 
  assign _2_8_io_x_px = _GEN_63[6]; 
  assign _2_8_io_x_pr = _GEN_63[5]; 
  assign _2_8_io_x_pal = _GEN_63[4];
  assign _2_8_io_x_paa = _GEN_63[3];
  assign _2_8_io_x_eff = _GEN_63[2];
  assign _2_8_io_x_c = _GEN_63[1];

  assign _2_9_io_x_ppn = superpage_entries_0_data_0[33:14];
  assign _2_9_io_x_u = superpage_entries_0_data_0[13]; 
  assign _2_9_io_x_ae = superpage_entries_0_data_0[11];
  assign _2_9_io_x_sw = superpage_entries_0_data_0[10];
  assign _2_9_io_x_sx = superpage_entries_0_data_0[9]; 
  assign _2_9_io_x_sr = superpage_entries_0_data_0[8]; 
  assign _2_9_io_x_pw = superpage_entries_0_data_0[7]; 
  assign _2_9_io_x_px = superpage_entries_0_data_0[6]; 
  assign _2_9_io_x_pr = superpage_entries_0_data_0[5]; 
  assign _2_9_io_x_pal = superpage_entries_0_data_0[4];
  assign _2_9_io_x_paa = superpage_entries_0_data_0[3];
  assign _2_9_io_x_eff = superpage_entries_0_data_0[2];
  assign _2_9_io_x_c = superpage_entries_0_data_0[1];
  assign _2_10_io_x_ppn = superpage_entries_1_data_0[33:14];
  assign _2_10_io_x_u = superpage_entries_1_data_0[13]; 
  assign _2_10_io_x_ae = superpage_entries_1_data_0[11];
  assign _2_10_io_x_sw = superpage_entries_1_data_0[10];
  assign _2_10_io_x_sx = superpage_entries_1_data_0[9]; 
  assign _2_10_io_x_sr = superpage_entries_1_data_0[8]; 
  assign _2_10_io_x_pw = superpage_entries_1_data_0[7]; 
  assign _2_10_io_x_px = superpage_entries_1_data_0[6]; 
  assign _2_10_io_x_pr = superpage_entries_1_data_0[5]; 
  assign _2_10_io_x_pal = superpage_entries_1_data_0[4];
  assign _2_10_io_x_paa = superpage_entries_1_data_0[3];
  assign _2_10_io_x_eff = superpage_entries_1_data_0[2];
  assign _2_10_io_x_c = superpage_entries_1_data_0[1];
  assign _2_11_io_x_ppn = superpage_entries_2_data_0[33:14];
  assign _2_11_io_x_u = superpage_entries_2_data_0[13]; 
  assign _2_11_io_x_ae = superpage_entries_2_data_0[11];
  assign _2_11_io_x_sw = superpage_entries_2_data_0[10];
  assign _2_11_io_x_sx = superpage_entries_2_data_0[9]; 
  assign _2_11_io_x_sr = superpage_entries_2_data_0[8]; 
  assign _2_11_io_x_pw = superpage_entries_2_data_0[7]; 
  assign _2_11_io_x_px = superpage_entries_2_data_0[6]; 
  assign _2_11_io_x_pr = superpage_entries_2_data_0[5]; 
  assign _2_11_io_x_pal = superpage_entries_2_data_0[4];
  assign _2_11_io_x_paa = superpage_entries_2_data_0[3];
  assign _2_11_io_x_eff = superpage_entries_2_data_0[2];
  assign _2_11_io_x_c = superpage_entries_2_data_0[1];
  assign _2_12_io_x_ppn = superpage_entries_3_data_0[33:14];
  assign _2_12_io_x_u = superpage_entries_3_data_0[13]; 
  assign _2_12_io_x_ae = superpage_entries_3_data_0[11];
  assign _2_12_io_x_sw = superpage_entries_3_data_0[10];
  assign _2_12_io_x_sx = superpage_entries_3_data_0[9]; 
  assign _2_12_io_x_sr = superpage_entries_3_data_0[8]; 
  assign _2_12_io_x_pw = superpage_entries_3_data_0[7]; 
  assign _2_12_io_x_px = superpage_entries_3_data_0[6]; 
  assign _2_12_io_x_pr = superpage_entries_3_data_0[5]; 
  assign _2_12_io_x_pal = superpage_entries_3_data_0[4];
  assign _2_12_io_x_paa = superpage_entries_3_data_0[3];
  assign _2_12_io_x_eff = superpage_entries_3_data_0[2];
  assign _2_12_io_x_c = superpage_entries_3_data_0[1];
  assign _2_13_io_x_ppn = special_entry_data_0[33:14];
  assign _2_13_io_x_u = special_entry_data_0[13]; 
  assign _2_13_io_x_ae = special_entry_data_0[11];
  assign _2_13_io_x_sw = special_entry_data_0[10];
  assign _2_13_io_x_sx = special_entry_data_0[9]; 
  assign _2_13_io_x_sr = special_entry_data_0[8]; 
  assign _2_13_io_x_pw = special_entry_data_0[7]; 
  assign _2_13_io_x_px = special_entry_data_0[6]; 
  assign _2_13_io_x_pr = special_entry_data_0[5]; 
  assign _2_13_io_x_pal = special_entry_data_0[4];
  assign _2_13_io_x_paa = special_entry_data_0[3];
  assign _2_13_io_x_eff = special_entry_data_0[2];
  assign _2_13_io_x_c = special_entry_data_0[1]; 

  assign _2_14_io_x_ppn = _GEN_35[33:14];
  assign _2_14_io_x_u = _GEN_35[13];
  assign _2_14_io_x_ae = _GEN_35[11];
  assign _2_14_io_x_sw = _GEN_35[10];
  assign _2_14_io_x_sx = _GEN_35[9];
  assign _2_14_io_x_sr = _GEN_35[8];
  assign _2_14_io_x_pw = _GEN_35[7];
  assign _2_14_io_x_px = _GEN_35[6];
  assign _2_14_io_x_pr = _GEN_35[5];
  assign _2_14_io_x_pal = _GEN_35[4];
  assign _2_14_io_x_paa = _GEN_35[3];
  assign _2_14_io_x_eff = _GEN_35[2];
  assign _2_14_io_x_c = _GEN_35[1];
  assign _2_15_io_x_ppn = _GEN_39[33:14];
  assign _2_15_io_x_u = _GEN_39[13];
  assign _2_15_io_x_ae = _GEN_39[11];
  assign _2_15_io_x_sw = _GEN_39[10];
  assign _2_15_io_x_sx = _GEN_39[9];
  assign _2_15_io_x_sr = _GEN_39[8];
  assign _2_15_io_x_pw = _GEN_39[7];
  assign _2_15_io_x_px = _GEN_39[6];
  assign _2_15_io_x_pr = _GEN_39[5];
  assign _2_15_io_x_pal = _GEN_39[4];
  assign _2_15_io_x_paa = _GEN_39[3];
  assign _2_15_io_x_eff = _GEN_39[2];
  assign _2_15_io_x_c = _GEN_39[1];
  assign _2_16_io_x_ppn = _GEN_43[33:14];
  assign _2_16_io_x_u = _GEN_43[13];
  assign _2_16_io_x_ae = _GEN_43[11];
  assign _2_16_io_x_sw = _GEN_43[10];
  assign _2_16_io_x_sx = _GEN_43[9];
  assign _2_16_io_x_sr = _GEN_43[8];
  assign _2_16_io_x_pw = _GEN_43[7];
  assign _2_16_io_x_px = _GEN_43[6];
  assign _2_16_io_x_pr = _GEN_43[5];
  assign _2_16_io_x_pal = _GEN_43[4];
  assign _2_16_io_x_paa = _GEN_43[3];
  assign _2_16_io_x_eff = _GEN_43[2];
  assign _2_16_io_x_c = _GEN_43[1];
  assign _2_17_io_x_ppn = _GEN_47[33:14];
  assign _2_17_io_x_u = _GEN_47[13];
  assign _2_17_io_x_ae = _GEN_47[11];
  assign _2_17_io_x_sw = _GEN_47[10];
  assign _2_17_io_x_sx = _GEN_47[9];
  assign _2_17_io_x_sr = _GEN_47[8];
  assign _2_17_io_x_pw = _GEN_47[7];
  assign _2_17_io_x_px = _GEN_47[6];
  assign _2_17_io_x_pr = _GEN_47[5];
  assign _2_17_io_x_pal = _GEN_47[4];
  assign _2_17_io_x_paa = _GEN_47[3];
  assign _2_17_io_x_eff = _GEN_47[2];
  assign _2_17_io_x_c = _GEN_47[1];
  assign _2_18_io_x_ppn = _GEN_51[33:14];
  assign _2_18_io_x_u = _GEN_51[13];
  assign _2_18_io_x_ae = _GEN_51[11];
  assign _2_18_io_x_sw = _GEN_51[10];
  assign _2_18_io_x_sx = _GEN_51[9];
  assign _2_18_io_x_sr = _GEN_51[8];
  assign _2_18_io_x_pw = _GEN_51[7];
  assign _2_18_io_x_px = _GEN_51[6];
  assign _2_18_io_x_pr = _GEN_51[5];
  assign _2_18_io_x_pal = _GEN_51[4];
  assign _2_18_io_x_paa = _GEN_51[3];
  assign _2_18_io_x_eff = _GEN_51[2];
  assign _2_18_io_x_c = _GEN_51[1];
  assign _2_19_io_x_ppn = _GEN_55[33:14];
  assign _2_19_io_x_u = _GEN_55[13];
  assign _2_19_io_x_ae = _GEN_55[11];
  assign _2_19_io_x_sw = _GEN_55[10];
  assign _2_19_io_x_sx = _GEN_55[9];
  assign _2_19_io_x_sr = _GEN_55[8];
  assign _2_19_io_x_pw = _GEN_55[7];
  assign _2_19_io_x_px = _GEN_55[6];
  assign _2_19_io_x_pr = _GEN_55[5];
  assign _2_19_io_x_pal = _GEN_55[4];
  assign _2_19_io_x_paa = _GEN_55[3];
  assign _2_19_io_x_eff = _GEN_55[2];
  assign _2_19_io_x_c = _GEN_55[1];
  assign _2_20_io_x_ppn = _GEN_59[33:14];
  assign _2_20_io_x_u = _GEN_59[13];
  assign _2_20_io_x_ae = _GEN_59[11];
  assign _2_20_io_x_sw = _GEN_59[10];
  assign _2_20_io_x_sx = _GEN_59[9];
  assign _2_20_io_x_sr = _GEN_59[8];
  assign _2_20_io_x_pw = _GEN_59[7];
  assign _2_20_io_x_px = _GEN_59[6];
  assign _2_20_io_x_pr = _GEN_59[5];
  assign _2_20_io_x_pal = _GEN_59[4];
  assign _2_20_io_x_paa = _GEN_59[3];
  assign _2_20_io_x_eff = _GEN_59[2];
  assign _2_20_io_x_c = _GEN_59[1];
  assign _2_21_io_x_ppn = _GEN_63[33:14];
  assign _2_21_io_x_u = _GEN_63[13];
  assign _2_21_io_x_ae = _GEN_63[11];
  assign _2_21_io_x_sw = _GEN_63[10];
  assign _2_21_io_x_sx = _GEN_63[9];
  assign _2_21_io_x_sr = _GEN_63[8];
  assign _2_21_io_x_pw = _GEN_63[7];
  assign _2_21_io_x_px = _GEN_63[6];
  assign _2_21_io_x_pr = _GEN_63[5]; 
  assign _2_21_io_x_pal = _GEN_63[4];
  assign _2_21_io_x_paa = _GEN_63[3];
  assign _2_21_io_x_eff = _GEN_63[2];
  assign _2_21_io_x_c = _GEN_63[1];

  assign _2_22_io_x_ppn = superpage_entries_0_data_0[33:14];
  assign _2_22_io_x_u = superpage_entries_0_data_0[13];
  assign _2_22_io_x_ae = superpage_entries_0_data_0[11];
  assign _2_22_io_x_sw = superpage_entries_0_data_0[10]; 
  assign _2_22_io_x_sx = superpage_entries_0_data_0[9];
  assign _2_22_io_x_sr = superpage_entries_0_data_0[8];
  assign _2_22_io_x_pw = superpage_entries_0_data_0[7];
  assign _2_22_io_x_px = superpage_entries_0_data_0[6];
  assign _2_22_io_x_pr = superpage_entries_0_data_0[5];
  assign _2_22_io_x_pal = superpage_entries_0_data_0[4];
  assign _2_22_io_x_paa = superpage_entries_0_data_0[3];
  assign _2_22_io_x_eff = superpage_entries_0_data_0[2];
  assign _2_22_io_x_c = superpage_entries_0_data_0[1];
  assign _2_23_io_x_ppn = superpage_entries_1_data_0[33:14];
  assign _2_23_io_x_u = superpage_entries_1_data_0[13];
  assign _2_23_io_x_ae = superpage_entries_1_data_0[11];
  assign _2_23_io_x_sw = superpage_entries_1_data_0[10];
  assign _2_23_io_x_sx = superpage_entries_1_data_0[9];
  assign _2_23_io_x_sr = superpage_entries_1_data_0[8];
  assign _2_23_io_x_pw = superpage_entries_1_data_0[7];
  assign _2_23_io_x_px = superpage_entries_1_data_0[6];
  assign _2_23_io_x_pr = superpage_entries_1_data_0[5];
  assign _2_23_io_x_pal = superpage_entries_1_data_0[4];
  assign _2_23_io_x_paa = superpage_entries_1_data_0[3];
  assign _2_23_io_x_eff = superpage_entries_1_data_0[2];
  assign _2_23_io_x_c = superpage_entries_1_data_0[1];
  assign _2_24_io_x_ppn = superpage_entries_2_data_0[33:14];
  assign _2_24_io_x_u = superpage_entries_2_data_0[13];
  assign _2_24_io_x_ae = superpage_entries_2_data_0[11];
  assign _2_24_io_x_sw = superpage_entries_2_data_0[10];
  assign _2_24_io_x_sx = superpage_entries_2_data_0[9];
  assign _2_24_io_x_sr = superpage_entries_2_data_0[8];
  assign _2_24_io_x_pw = superpage_entries_2_data_0[7];
  assign _2_24_io_x_px = superpage_entries_2_data_0[6]; 
  assign _2_24_io_x_pr = superpage_entries_2_data_0[5];
  assign _2_24_io_x_pal = superpage_entries_2_data_0[4];
  assign _2_24_io_x_paa = superpage_entries_2_data_0[3]; 
  assign _2_24_io_x_eff = superpage_entries_2_data_0[2];
  assign _2_24_io_x_c = superpage_entries_2_data_0[1];
  assign _2_25_io_x_ppn = superpage_entries_3_data_0[33:14];
  assign _2_25_io_x_u = superpage_entries_3_data_0[13];
  assign _2_25_io_x_ae = superpage_entries_3_data_0[11];
  assign _2_25_io_x_sw = superpage_entries_3_data_0[10];
  assign _2_25_io_x_sx = superpage_entries_3_data_0[9];
  assign _2_25_io_x_sr = superpage_entries_3_data_0[8];
  assign _2_25_io_x_pw = superpage_entries_3_data_0[7];
  assign _2_25_io_x_px = superpage_entries_3_data_0[6];
  assign _2_25_io_x_pr = superpage_entries_3_data_0[5];
  assign _2_25_io_x_pal = superpage_entries_3_data_0[4];
  assign _2_25_io_x_paa = superpage_entries_3_data_0[3];
  assign _2_25_io_x_eff = superpage_entries_3_data_0[2];
  assign _2_25_io_x_c = superpage_entries_3_data_0[1];
  assign _2_26_io_x_ppn = special_entry_data_0[33:14];
  assign _2_26_io_x_u = special_entry_data_0[13];
  assign _2_26_io_x_ae = special_entry_data_0[11];
  assign _2_26_io_x_sw = special_entry_data_0[10];
  assign _2_26_io_x_sx = special_entry_data_0[9];
  assign _2_26_io_x_sr = special_entry_data_0[8];
  assign _2_26_io_x_pw = special_entry_data_0[7];
  assign _2_26_io_x_px = special_entry_data_0[6];
  assign _2_26_io_x_pr = special_entry_data_0[5]; 
  assign _2_26_io_x_pal = special_entry_data_0[4];
  assign _2_26_io_x_paa = special_entry_data_0[3];
  assign _2_26_io_x_eff = special_entry_data_0[2];
  assign _2_26_io_x_c = special_entry_data_0[1];

  assign _2_27_io_x_ppn = _GEN_35[33:14];
  assign _2_27_io_x_u = _GEN_35[13];
  assign _2_27_io_x_ae = _GEN_35[11];
  assign _2_27_io_x_sw = _GEN_35[10];
  assign _2_27_io_x_sx = _GEN_35[9];
  assign _2_27_io_x_sr = _GEN_35[8];
  assign _2_27_io_x_pw = _GEN_35[7];
  assign _2_27_io_x_px = _GEN_35[6];
  assign _2_27_io_x_pr = _GEN_35[5];
  assign _2_27_io_x_pal = _GEN_35[4];
  assign _2_27_io_x_paa = _GEN_35[3];
  assign _2_27_io_x_eff = _GEN_35[2];
  assign _2_27_io_x_c = _GEN_35[1];
  assign _2_28_io_x_ppn = _GEN_39[33:14];
  assign _2_28_io_x_u = _GEN_39[13];
  assign _2_28_io_x_ae = _GEN_39[11];
  assign _2_28_io_x_sw = _GEN_39[10];
  assign _2_28_io_x_sx = _GEN_39[9];
  assign _2_28_io_x_sr = _GEN_39[8];
  assign _2_28_io_x_pw = _GEN_39[7];
  assign _2_28_io_x_px = _GEN_39[6];
  assign _2_28_io_x_pr = _GEN_39[5];
  assign _2_28_io_x_pal = _GEN_39[4];
  assign _2_28_io_x_paa = _GEN_39[3];
  assign _2_28_io_x_eff = _GEN_39[2];
  assign _2_28_io_x_c = _GEN_39[1]; 
  assign _2_29_io_x_ppn = _GEN_43[33:14];
  assign _2_29_io_x_u = _GEN_43[13];
  assign _2_29_io_x_ae = _GEN_43[11];
  assign _2_29_io_x_sw = _GEN_43[10];
  assign _2_29_io_x_sx = _GEN_43[9];
  assign _2_29_io_x_sr = _GEN_43[8];
  assign _2_29_io_x_pw = _GEN_43[7];
  assign _2_29_io_x_px = _GEN_43[6];
  assign _2_29_io_x_pr = _GEN_43[5];
  assign _2_29_io_x_pal = _GEN_43[4];
  assign _2_29_io_x_paa = _GEN_43[3];
  assign _2_29_io_x_eff = _GEN_43[2];
  assign _2_29_io_x_c = _GEN_43[1];
  assign _2_30_io_x_ppn = _GEN_47[33:14];
  assign _2_30_io_x_u = _GEN_47[13];
  assign _2_30_io_x_ae = _GEN_47[11];
  assign _2_30_io_x_sw = _GEN_47[10];
  assign _2_30_io_x_sx = _GEN_47[9];
  assign _2_30_io_x_sr = _GEN_47[8];
  assign _2_30_io_x_pw = _GEN_47[7];
  assign _2_30_io_x_px = _GEN_47[6];
  assign _2_30_io_x_pr = _GEN_47[5];
  assign _2_30_io_x_pal = _GEN_47[4];
  assign _2_30_io_x_paa = _GEN_47[3];
  assign _2_30_io_x_eff = _GEN_47[2];
  assign _2_30_io_x_c = _GEN_47[1];
  assign _2_31_io_x_ppn = _GEN_51[33:14];
  assign _2_31_io_x_u = _GEN_51[13];
  assign _2_31_io_x_ae = _GEN_51[11];
  assign _2_31_io_x_sw = _GEN_51[10];
  assign _2_31_io_x_sx = _GEN_51[9];
  assign _2_31_io_x_sr = _GEN_51[8];
  assign _2_31_io_x_pw = _GEN_51[7];
  assign _2_31_io_x_px = _GEN_51[6];
  assign _2_31_io_x_pr = _GEN_51[5];
  assign _2_31_io_x_pal = _GEN_51[4];
  assign _2_31_io_x_paa = _GEN_51[3];
  assign _2_31_io_x_eff = _GEN_51[2];
  assign _2_31_io_x_c = _GEN_51[1];
  assign _2_32_io_x_ppn = _GEN_55[33:14];
  assign _2_32_io_x_u = _GEN_55[13];
  assign _2_32_io_x_ae = _GEN_55[11];
  assign _2_32_io_x_sw = _GEN_55[10];
  assign _2_32_io_x_sx = _GEN_55[9];
  assign _2_32_io_x_sr = _GEN_55[8];
  assign _2_32_io_x_pw = _GEN_55[7];
  assign _2_32_io_x_px = _GEN_55[6];
  assign _2_32_io_x_pr = _GEN_55[5];
  assign _2_32_io_x_pal = _GEN_55[4];
  assign _2_32_io_x_paa = _GEN_55[3];
  assign _2_32_io_x_eff = _GEN_55[2];
  assign _2_32_io_x_c = _GEN_55[1];
  assign _2_33_io_x_ppn = _GEN_59[33:14];
  assign _2_33_io_x_u = _GEN_59[13];
  assign _2_33_io_x_ae = _GEN_59[11];
  assign _2_33_io_x_sw = _GEN_59[10];
  assign _2_33_io_x_sx = _GEN_59[9];
  assign _2_33_io_x_sr = _GEN_59[8];
  assign _2_33_io_x_pw = _GEN_59[7];
  assign _2_33_io_x_px = _GEN_59[6];
  assign _2_33_io_x_pr = _GEN_59[5];
  assign _2_33_io_x_pal = _GEN_59[4];
  assign _2_33_io_x_paa = _GEN_59[3];
  assign _2_33_io_x_eff = _GEN_59[2];
  assign _2_33_io_x_c = _GEN_59[1];
  assign _2_34_io_x_ppn = _GEN_63[33:14];
  assign _2_34_io_x_u = _GEN_63[13];
  assign _2_34_io_x_ae = _GEN_63[11];
  assign _2_34_io_x_sw = _GEN_63[10];
  assign _2_34_io_x_sx = _GEN_63[9];
  assign _2_34_io_x_sr = _GEN_63[8];
  assign _2_34_io_x_pw = _GEN_63[7];
  assign _2_34_io_x_px = _GEN_63[6];
  assign _2_34_io_x_pr = _GEN_63[5];
  assign _2_34_io_x_pal = _GEN_63[4];
  assign _2_34_io_x_paa = _GEN_63[3];
  assign _2_34_io_x_eff = _GEN_63[2];
  assign _2_34_io_x_c = _GEN_63[1];

  assign _2_35_io_x_ppn = superpage_entries_0_data_0[33:14];
  assign _2_35_io_x_u = superpage_entries_0_data_0[13];
  assign _2_35_io_x_ae = superpage_entries_0_data_0[11];
  assign _2_35_io_x_sw = superpage_entries_0_data_0[10];
  assign _2_35_io_x_sx = superpage_entries_0_data_0[9];
  assign _2_35_io_x_sr = superpage_entries_0_data_0[8];
  assign _2_35_io_x_pw = superpage_entries_0_data_0[7];
  assign _2_35_io_x_px = superpage_entries_0_data_0[6];
  assign _2_35_io_x_pr = superpage_entries_0_data_0[5];
  assign _2_35_io_x_pal = superpage_entries_0_data_0[4];
  assign _2_35_io_x_paa = superpage_entries_0_data_0[3];
  assign _2_35_io_x_eff = superpage_entries_0_data_0[2];
  assign _2_35_io_x_c = superpage_entries_0_data_0[1];
  assign _2_36_io_x_ppn = superpage_entries_1_data_0[33:14];
  assign _2_36_io_x_u = superpage_entries_1_data_0[13];
  assign _2_36_io_x_ae = superpage_entries_1_data_0[11];
  assign _2_36_io_x_sw = superpage_entries_1_data_0[10];
  assign _2_36_io_x_sx = superpage_entries_1_data_0[9];
  assign _2_36_io_x_sr = superpage_entries_1_data_0[8];
  assign _2_36_io_x_pw = superpage_entries_1_data_0[7];
  assign _2_36_io_x_px = superpage_entries_1_data_0[6];
  assign _2_36_io_x_pr = superpage_entries_1_data_0[5];
  assign _2_36_io_x_pal = superpage_entries_1_data_0[4];
  assign _2_36_io_x_paa = superpage_entries_1_data_0[3];
  assign _2_36_io_x_eff = superpage_entries_1_data_0[2];
  assign _2_36_io_x_c = superpage_entries_1_data_0[1];
  assign _2_37_io_x_ppn = superpage_entries_2_data_0[33:14];
  assign _2_37_io_x_u = superpage_entries_2_data_0[13];
  assign _2_37_io_x_ae = superpage_entries_2_data_0[11];
  assign _2_37_io_x_sw = superpage_entries_2_data_0[10];
  assign _2_37_io_x_sx = superpage_entries_2_data_0[9];
  assign _2_37_io_x_sr = superpage_entries_2_data_0[8];
  assign _2_37_io_x_pw = superpage_entries_2_data_0[7];
  assign _2_37_io_x_px = superpage_entries_2_data_0[6];
  assign _2_37_io_x_pr = superpage_entries_2_data_0[5];
  assign _2_37_io_x_pal = superpage_entries_2_data_0[4];
  assign _2_37_io_x_paa = superpage_entries_2_data_0[3];
  assign _2_37_io_x_eff = superpage_entries_2_data_0[2];
  assign _2_37_io_x_c = superpage_entries_2_data_0[1];
  assign _2_38_io_x_ppn = superpage_entries_3_data_0[33:14];
  assign _2_38_io_x_u = superpage_entries_3_data_0[13];
  assign _2_38_io_x_ae = superpage_entries_3_data_0[11];
  assign _2_38_io_x_sw = superpage_entries_3_data_0[10];
  assign _2_38_io_x_sx = superpage_entries_3_data_0[9];
  assign _2_38_io_x_sr = superpage_entries_3_data_0[8];
  assign _2_38_io_x_pw = superpage_entries_3_data_0[7];
  assign _2_38_io_x_px = superpage_entries_3_data_0[6];
  assign _2_38_io_x_pr = superpage_entries_3_data_0[5]; 
  assign _2_38_io_x_pal = superpage_entries_3_data_0[4];
  assign _2_38_io_x_paa = superpage_entries_3_data_0[3];
  assign _2_38_io_x_eff = superpage_entries_3_data_0[2];
  assign _2_38_io_x_c = superpage_entries_3_data_0[1];
//Passed

  wire _T_893 = io_ptw_resp_valid & !invalidate_refill;
  wire _T_900 = io_ptw_resp_bits_pte_v & (io_ptw_resp_bits_pte_r | (io_ptw_resp_bits_pte_x & !io_ptw_resp_bits_pte_w)) & io_ptw_resp_bits_pte_a;
  wire _T_915 = io_ptw_resp_bits_homogeneous == 1'h0;
  wire [33:0] _T_931 = {refill_ppn
		,io_ptw_resp_bits_pte_u
		,(io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v)
		,io_ptw_resp_bits_ae
		,(_T_900 & io_ptw_resp_bits_pte_w & io_ptw_resp_bits_pte_d)
		,(_T_900 & io_ptw_resp_bits_pte_x)
		,(_T_900 & io_ptw_resp_bits_pte_r)
		,prot_w
		,prot_x,prot_r,prot_al,prot_al,prot_eff,cacheable,1'h0}; 
  wire _T_932 = io_ptw_resp_bits_level < 1'h1;
  wire [2:0] _T_993 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; 
  wire _T_994 = _T_993 == 3'h0;
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & !(_T_932) & _T_994) begin
		sectored_entries_0_tag <= r_refill_tag;
		if (2'h0 == r_refill_tag[1:0]) begin
			sectored_entries_0_data_0 <= _T_931;
		end
		if (2'h1 == r_refill_tag[1:0]) begin
			sectored_entries_0_data_1 <= _T_931;
		end
		if (2'h2 == r_refill_tag[1:0]) begin
			sectored_entries_0_data_2 <= _T_931;
		end
		if (2'h3 == r_refill_tag[1:0]) begin
			sectored_entries_0_data_3 <= _T_931;
		end
	end
end

  wire _T_2258 = _T_380[19:10] == 10'h0;
  wire _T_3589 = multipleHits | reset;
  wire _GEN_950 = 2'h0 == r_refill_tag[1:0];
  wire _T_995 = r_sectored_hit == 1'h0;
  wire _GEN_84 = _GEN_950 
		| (_T_995 ? 1'h0 : sectored_entries_0_valid_0);
  wire _GEN_472 = !_T_893 ? sectored_entries_0_valid_0
			: _T_915 ? sectored_entries_0_valid_0 
			: _T_932 ? sectored_entries_0_valid_0 
			: _T_994 ? _GEN_84 
			: sectored_entries_0_valid_0;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_0_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2258 & sectored_entries_0_data_0[0]) begin
				    sectored_entries_0_valid_0 <= 1'h0;
				end else begin
					if (_T_382 & (2'h0 == _T_477)) begin
						sectored_entries_0_valid_0 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_994) begin
							sectored_entries_0_valid_0 <= _GEN_84;
						end
					end
				end
			end else begin
				sectored_entries_0_valid_0 <= io_sfence_bits_rs2 & (!sectored_entries_0_data_0[12] ? 1'h0 : _GEN_472);
			end
		end else begin
			sectored_entries_0_valid_0 <= _GEN_472;
		end
	end
end
// Passed
  wire _GEN_951 = 2'h1 == r_refill_tag[1:0];
  wire _GEN_85 = _GEN_951 
		| (_T_995 ? 1'h0 : sectored_entries_0_valid_1);
  wire _GEN_473 = !_T_893 ? sectored_entries_0_valid_1
			: _T_915 ? sectored_entries_0_valid_1 
			: _T_932 ? sectored_entries_0_valid_1 
			: _T_994 ? _GEN_85 
			: sectored_entries_0_valid_1;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_0_valid_1 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2258 & sectored_entries_0_data_1[0]) begin
				    sectored_entries_0_valid_1 <= 1'h0;
				end else begin
					if (_T_382 & (2'h1 == _T_477)) begin
						sectored_entries_0_valid_1 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_994) begin
							sectored_entries_0_valid_1 <= _GEN_85;
						end
					end
				end
			end else begin
				sectored_entries_0_valid_1 <= io_sfence_bits_rs2 & (!sectored_entries_0_data_1[12] ? 1'h0 : _GEN_473);
			end
		end else begin
			sectored_entries_0_valid_1 <= _GEN_473;
		end
	end
end
// Passed 
  wire _GEN_952 = 2'h2 == r_refill_tag[1:0];
  wire _GEN_86 = _GEN_952 
  		| (_T_995 ? 1'h0 : sectored_entries_0_valid_2);
  wire _GEN_474 = !_T_893 ? sectored_entries_0_valid_2
			: _T_915 ? sectored_entries_0_valid_2 
			: _T_932 ? sectored_entries_0_valid_2 
			: _T_994 ? _GEN_86 
			: sectored_entries_0_valid_2;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_0_valid_2 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2258 & sectored_entries_0_data_2[0]) begin
				    sectored_entries_0_valid_2 <= 1'h0;
				end else begin
					if (_T_382 & (2'h2 == _T_477)) begin
						sectored_entries_0_valid_2 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_994) begin
							sectored_entries_0_valid_2 <= _GEN_86;
						end
					end
				end
			end else begin
				sectored_entries_0_valid_2 <= io_sfence_bits_rs2 & (!sectored_entries_0_data_2[12] ? 1'h0 : _GEN_474);
			end
		end else begin
			sectored_entries_0_valid_2 <= _GEN_474;
		end
	end
end

  wire _GEN_953 = 2'h3 == r_refill_tag[1:0];
  wire _GEN_87 = _GEN_953 
		| (_T_995 ? 1'h0 : sectored_entries_0_valid_3);
  wire _GEN_475 = !_T_893 ? sectored_entries_0_valid_3
			: _T_915 ? sectored_entries_0_valid_3 
			: _T_932 ? sectored_entries_0_valid_3 
			: _T_994 ? _GEN_87 
			: sectored_entries_0_valid_3;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_0_valid_3 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2258 & sectored_entries_0_data_3[0]) begin
				    sectored_entries_0_valid_3 <= 1'h0;
				end else begin
					if (_T_382 & (2'h3 == _T_477)) begin
						sectored_entries_0_valid_3 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_994) begin
							sectored_entries_0_valid_3 <= _GEN_87;
						end
					end
				end
			end else begin
				sectored_entries_0_valid_3 <= io_sfence_bits_rs2 & (!sectored_entries_0_data_3[12] ? 1'h0 : _GEN_475);
			end
		end else begin
			sectored_entries_0_valid_3 <= _GEN_475;
		end
	end
end
// Passed
  wire _T_1011 = _T_993 == 3'h1;
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & !(_T_932) & _T_1011) begin
		sectored_entries_1_tag <= r_refill_tag;
		if (2'h0 == r_refill_tag[1:0]) begin
			sectored_entries_1_data_0 <= _T_931;
		end
		if (2'h1 == r_refill_tag[1:0]) begin
			sectored_entries_1_data_1 <= _T_931;
		end
		if (2'h2 == r_refill_tag[1:0]) begin
			sectored_entries_1_data_2 <= _T_931;
		end
		if (2'h3 == r_refill_tag[1:0]) begin
			sectored_entries_1_data_3 <= _T_931;
		end
	end
end

  wire _T_2405 = _T_386[19:10] == 10'h0;
  wire _GEN_106 = _GEN_950 
		| (_T_995 ? 1'h0 : sectored_entries_1_valid_0);
  wire _GEN_482 = !_T_893 ? sectored_entries_1_valid_0
			: _T_915 ? sectored_entries_1_valid_0 
			: _T_932 ? sectored_entries_1_valid_0 
			: _T_1011 ? _GEN_106 
			: sectored_entries_1_valid_0;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_1_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2405 & sectored_entries_1_data_0[0]) begin
				    sectored_entries_1_valid_0 <= 1'h0;
				end else begin
					if (_T_388 & (2'h0 == _T_477)) begin
						sectored_entries_1_valid_0 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1011) begin
							sectored_entries_1_valid_0 <= _GEN_106;
						end
					end
				end
			end else begin
				sectored_entries_1_valid_0 <= io_sfence_bits_rs2 & (!sectored_entries_1_data_0[12] ? 1'h0 : _GEN_482);
			end
		end else begin
			sectored_entries_1_valid_0 <= _GEN_482;
		end
	end
end

  wire _GEN_107 = _GEN_951 
		| (_T_995 ? 1'h0 : sectored_entries_1_valid_1);
  wire _GEN_483 = !_T_893 ? sectored_entries_1_valid_1
			: _T_915 ? sectored_entries_1_valid_1 
			: _T_932 ? sectored_entries_1_valid_1 
			: _T_1011 ? _GEN_107 
			: sectored_entries_1_valid_1;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_1_valid_1 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2405 & sectored_entries_1_data_1[0]) begin
				    sectored_entries_1_valid_1 <= 1'h0;
				end else begin
					if (_T_388 & (2'h0 == _T_477)) begin
						sectored_entries_1_valid_1 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1011) begin
							sectored_entries_1_valid_1 <= _GEN_107;
						end
					end
				end
			end else begin
				sectored_entries_1_valid_1 <= io_sfence_bits_rs2 & (!sectored_entries_1_data_1[12] ? 1'h0 : _GEN_483);
			end
		end else begin
			sectored_entries_1_valid_1 <= _GEN_483;
		end
	end
end

  wire _GEN_108 = _GEN_952 
		| (_T_995 ? 1'h0 : sectored_entries_1_valid_2);
  wire _GEN_484 = !_T_893 ? sectored_entries_1_valid_2
			: _T_915 ? sectored_entries_1_valid_2 
			: _T_932 ? sectored_entries_1_valid_2 
			: _T_1011 ? _GEN_108 
			: sectored_entries_1_valid_2;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_1_valid_2 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2405 & sectored_entries_1_data_2[0]) begin
				    sectored_entries_1_valid_2 <= 1'h0;
				end else begin
					if (_T_388 & (2'h0 == _T_477)) begin
						sectored_entries_1_valid_2 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1011) begin
							sectored_entries_1_valid_2 <= _GEN_108;
						end
					end
				end
			end else begin
				sectored_entries_1_valid_2 <= io_sfence_bits_rs2 & (!sectored_entries_1_data_2[12] ? 1'h0 : _GEN_484);
			end
		end else begin
			sectored_entries_1_valid_2 <= _GEN_484;
		end
	end
end

  wire _GEN_109 = _GEN_953 
		| (_T_995 ? 1'h0 : sectored_entries_1_valid_3);
  wire _GEN_485 = !_T_893 ? sectored_entries_1_valid_3
			: _T_915 ? sectored_entries_1_valid_3 
			: _T_932 ? sectored_entries_1_valid_3 
			: _T_1011 ? _GEN_109 
			: sectored_entries_1_valid_3;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_1_valid_3 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2405 & sectored_entries_1_data_3[0]) begin
				    sectored_entries_1_valid_3 <= 1'h0;
				end else begin
					if (_T_388 & (2'h0 == _T_477)) begin
						sectored_entries_1_valid_3 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1011) begin
							sectored_entries_1_valid_3 <= _GEN_109;
						end
					end
				end
			end else begin
				sectored_entries_1_valid_3 <= io_sfence_bits_rs2 & (!sectored_entries_1_data_3[12] ? 1'h0 : _GEN_485);
			end
		end else begin
			sectored_entries_1_valid_3 <= _GEN_485;
		end
	end
end

  wire _T_1028 = _T_993 == 3'h2;
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & !(_T_932) & _T_1028) begin
		sectored_entries_2_tag <= r_refill_tag;
		if (2'h0 == r_refill_tag[1:0]) begin
			sectored_entries_2_data_0 <= _T_931;
		end
		if (2'h1 == r_refill_tag[1:0]) begin
			sectored_entries_2_data_1 <= _T_931;
		end
		if (2'h2 == r_refill_tag[1:0]) begin
			sectored_entries_2_data_2 <= _T_931;
		end
		if (2'h3 == r_refill_tag[1:0]) begin
			sectored_entries_2_data_3 <= _T_931;
		end
	end
end

  wire _T_2552 = _T_392[19:10] == 10'h0;
  wire _GEN_128 = _GEN_950 
		| (_T_995 ? 1'h0 : sectored_entries_2_valid_0);
  wire _GEN_492 = !_T_893 ? sectored_entries_2_valid_0
			: _T_915 ? sectored_entries_2_valid_0 
			: _T_932 ? sectored_entries_2_valid_0 
			: _T_1028 ? _GEN_128 
			: sectored_entries_2_valid_0;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_2_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2552 & sectored_entries_2_data_0[0]) begin
				    sectored_entries_2_valid_0 <= 1'h0;
				end else begin
					if (_T_394 & (2'h0 == _T_477)) begin
						sectored_entries_2_valid_0 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1028) begin
							sectored_entries_2_valid_0 <= _GEN_128;
						end
					end
				end
			end else begin
				sectored_entries_2_valid_0 <= io_sfence_bits_rs2 & (!sectored_entries_2_data_0[12] ? 1'h0 : _GEN_492);
			end
		end else begin
			sectored_entries_2_valid_0 <= _GEN_492;
		end
	end
end

  wire _GEN_129 = _GEN_951 
		| (_T_995 ? 1'h0 : sectored_entries_2_valid_1);
  wire _GEN_493 = !_T_893 ? sectored_entries_2_valid_1
			: _T_915 ? sectored_entries_2_valid_1 
			: _T_932 ? sectored_entries_2_valid_1 
			: _T_1028 ? _GEN_129 
			: sectored_entries_2_valid_1;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_2_valid_1 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2552 & sectored_entries_2_data_1[0]) begin
				    sectored_entries_2_valid_1 <= 1'h0;
				end else begin
					if (_T_394 & (2'h0 == _T_477)) begin
						sectored_entries_2_valid_1 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1028) begin
							sectored_entries_2_valid_1 <= _GEN_129;
						end
					end
				end
			end else begin
				sectored_entries_2_valid_1 <= io_sfence_bits_rs2 & (!sectored_entries_2_data_1[12] ? 1'h0 : _GEN_493);
			end
		end else begin
			sectored_entries_2_valid_1 <= _GEN_493;
		end
	end
end

  wire _GEN_130 = _GEN_952 
		| (_T_995 ? 1'h0 : sectored_entries_2_valid_2);
  wire _GEN_494 = !_T_893 ? sectored_entries_2_valid_2
			: _T_915 ? sectored_entries_2_valid_2 
			: _T_932 ? sectored_entries_2_valid_2 
			: _T_1028 ? _GEN_130 
			: sectored_entries_2_valid_2;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_2_valid_2 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2552 & sectored_entries_2_data_2[0]) begin
				    sectored_entries_2_valid_2 <= 1'h0;
				end else begin
					if (_T_394 & (2'h0 == _T_477)) begin
						sectored_entries_2_valid_2 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1028) begin
							sectored_entries_2_valid_2 <= _GEN_130;
						end
					end
				end
			end else begin
				sectored_entries_2_valid_2 <= io_sfence_bits_rs2 & (!sectored_entries_2_data_2[12] ? 1'h0 : _GEN_494);
			end
		end else begin
			sectored_entries_2_valid_2 <= _GEN_494;
		end
	end
end

  wire _GEN_131 = _GEN_953 
		| (_T_995 ? 1'h0 : sectored_entries_2_valid_3);
  wire _GEN_495 = !_T_893 ? sectored_entries_2_valid_3
			: _T_915 ? sectored_entries_2_valid_3 
			: _T_932 ? sectored_entries_2_valid_3 
			: _T_1028 ? _GEN_131 
			: sectored_entries_2_valid_3;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_2_valid_3 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2552 & sectored_entries_2_data_3[0]) begin
				    sectored_entries_2_valid_3 <= 1'h0;
				end else begin
					if (_T_394 & (2'h0 == _T_477)) begin
						sectored_entries_2_valid_3 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1028) begin
							sectored_entries_2_valid_3 <= _GEN_131;
						end
					end
				end
			end else begin
				sectored_entries_2_valid_3 <= io_sfence_bits_rs2 & (!sectored_entries_2_data_3[12] ? 1'h0 : _GEN_495);
			end
		end else begin
			sectored_entries_2_valid_3 <= _GEN_495;
		end
	end
end
// Passed
  wire _T_1045 = _T_993 == 3'h3;
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & !(_T_932) & _T_1045) begin
		sectored_entries_3_tag <= r_refill_tag;
		if (2'h0 == r_refill_tag[1:0]) begin
			sectored_entries_3_data_0 <= _T_931;
		end
		if (2'h1 == r_refill_tag[1:0]) begin
			sectored_entries_3_data_1 <= _T_931;
		end
		if (2'h2 == r_refill_tag[1:0]) begin
			sectored_entries_3_data_2 <= _T_931;
		end
		if (2'h3 == r_refill_tag[1:0]) begin
			sectored_entries_3_data_3 <= _T_931;
		end
	end
end

  wire _T_2699 = _T_398[19:10] == 10'h0;
  wire _GEN_150 = _GEN_950 
		| (_T_995 ? 1'h0 : sectored_entries_3_valid_0);
  wire _GEN_502 = !_T_893 ? sectored_entries_3_valid_0
			: _T_915 ? sectored_entries_3_valid_0 
			: _T_932 ? sectored_entries_3_valid_0 
			: _T_1045 ? _GEN_150 
			: sectored_entries_3_valid_0;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_3_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2699 & sectored_entries_3_data_0[0]) begin
				    sectored_entries_3_valid_0 <= 1'h0;
				end else begin
					if (_T_400 & (2'h0 == _T_477)) begin
						sectored_entries_3_valid_0 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1045) begin
							sectored_entries_3_valid_0 <= _GEN_150;
						end
					end
				end
			end else begin
				sectored_entries_3_valid_0 <= io_sfence_bits_rs2 & (!sectored_entries_3_data_0[12] ? 1'h0 : _GEN_502);
			end
		end else begin
			sectored_entries_3_valid_0 <= _GEN_502;
		end
	end
end

  wire _GEN_151 = _GEN_951 
		| (_T_995 ? 1'h0 : sectored_entries_3_valid_1);
  wire _GEN_503 = !_T_893 ? sectored_entries_3_valid_1
			: _T_915 ? sectored_entries_3_valid_1 
			: _T_932 ? sectored_entries_3_valid_1 
			: _T_1045 ? _GEN_151 
			: sectored_entries_3_valid_1;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_3_valid_1 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2699 & sectored_entries_3_data_1[0]) begin
				    sectored_entries_3_valid_1 <= 1'h0;
				end else begin
					if (_T_400 & (2'h0 == _T_477)) begin
						sectored_entries_3_valid_1 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1045) begin
							sectored_entries_3_valid_1 <= _GEN_151;
						end
					end
				end
			end else begin
				sectored_entries_3_valid_1 <= io_sfence_bits_rs2 & (!sectored_entries_3_data_1[12] ? 1'h0 : _GEN_503);
			end
		end else begin
			sectored_entries_3_valid_1 <= _GEN_503;
		end
	end
end

  wire _GEN_152 = _GEN_952 
		| (_T_995 ? 1'h0 : sectored_entries_3_valid_2);
  wire _GEN_504 = !_T_893 ? sectored_entries_3_valid_2
			: _T_915 ? sectored_entries_3_valid_2 
			: _T_932 ? sectored_entries_3_valid_2 
			: _T_1045 ? _GEN_152 
			: sectored_entries_3_valid_2;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_3_valid_2 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2699 & sectored_entries_3_data_2[0]) begin
				    sectored_entries_3_valid_2 <= 1'h0;
				end else begin
					if (_T_400 & (2'h0 == _T_477)) begin
						sectored_entries_3_valid_2 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1045) begin
							sectored_entries_3_valid_2 <= _GEN_152;
						end
					end
				end
			end else begin
				sectored_entries_3_valid_2 <= io_sfence_bits_rs2 & (!sectored_entries_3_data_2[12] ? 1'h0 : _GEN_504);
			end
		end else begin
			sectored_entries_3_valid_2 <= _GEN_504;
		end
	end
end

  wire _GEN_153 = _GEN_953 
		| (_T_995 ? 1'h0 : sectored_entries_3_valid_3);
  wire _GEN_505 = !_T_893 ? sectored_entries_3_valid_3
			: _T_915 ? sectored_entries_3_valid_3 
			: _T_932 ? sectored_entries_3_valid_3 
			: _T_1045 ? _GEN_153 
			: sectored_entries_3_valid_3;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_3_valid_3 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2699 & sectored_entries_3_data_3[0]) begin
				    sectored_entries_3_valid_3 <= 1'h0;
				end else begin
					if (_T_400 & (2'h0 == _T_477)) begin
						sectored_entries_3_valid_3 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1045) begin
							sectored_entries_3_valid_3 <= _GEN_153;
						end
					end
				end
			end else begin
				sectored_entries_3_valid_3 <= io_sfence_bits_rs2 & (!sectored_entries_3_data_3[12] ? 1'h0 : _GEN_505);
			end
		end else begin
			sectored_entries_3_valid_3 <= _GEN_505;
		end
	end
end

  wire _T_1062 = _T_993 == 3'h4;
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & !(_T_932) & _T_1062) begin
		sectored_entries_4_tag <= r_refill_tag;
		if (2'h0 == r_refill_tag[1:0]) begin
			sectored_entries_4_data_0 <= _T_931;
		end
		if (2'h1 == r_refill_tag[1:0]) begin
			sectored_entries_4_data_1 <= _T_931;
		end
		if (2'h2 == r_refill_tag[1:0]) begin
			sectored_entries_4_data_2 <= _T_931;
		end
		if (2'h3 == r_refill_tag[1:0]) begin
			sectored_entries_4_data_3 <= _T_931;
		end
	end
end

  wire _T_2846 = _T_404[19:10] == 10'h0;
  wire _GEN_172 = _GEN_950 
		| (_T_995 ? 1'h0 : sectored_entries_4_valid_0);
  wire _GEN_512 = !_T_893 ? sectored_entries_4_valid_0
			: _T_915 ? sectored_entries_4_valid_0 
			: _T_932 ? sectored_entries_4_valid_0 
			: _T_1062 ? _GEN_172 
			: sectored_entries_4_valid_0;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_4_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2846 & sectored_entries_4_data_0[0]) begin
				    sectored_entries_4_valid_0 <= 1'h0;
				end else begin
					if (_T_406 & (2'h0 == _T_477)) begin
						sectored_entries_4_valid_0 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1062) begin
							sectored_entries_4_valid_0 <= _GEN_172;
						end
					end
				end
			end else begin
				sectored_entries_4_valid_0 <= io_sfence_bits_rs2 & (!sectored_entries_4_data_0[12] ? 1'h0 : _GEN_512);
			end
		end else begin
			sectored_entries_4_valid_0 <= _GEN_512;
		end
	end
end

  wire _GEN_173 = _GEN_951 
		| (_T_995 ? 1'h0 : sectored_entries_4_valid_1);
  wire _GEN_513 = !_T_893 ? sectored_entries_4_valid_1
			: _T_915 ? sectored_entries_4_valid_1 
			: _T_932 ? sectored_entries_4_valid_1 
			: _T_1062 ? _GEN_173 
			: sectored_entries_4_valid_1;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_4_valid_1 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2846 & sectored_entries_4_data_1[0]) begin
				    sectored_entries_4_valid_1 <= 1'h0;
				end else begin
					if (_T_406 & (2'h0 == _T_477)) begin
						sectored_entries_4_valid_1 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1062) begin
							sectored_entries_4_valid_1 <= _GEN_173;
						end
					end
				end
			end else begin
				sectored_entries_4_valid_1 <= io_sfence_bits_rs2 & (!sectored_entries_4_data_1[12] ? 1'h0 : _GEN_513);
			end
		end else begin
			sectored_entries_4_valid_1 <= _GEN_513;
		end
	end
end

  wire _GEN_174 = _GEN_952 
		| (_T_995 ? 1'h0 : sectored_entries_4_valid_2);
  wire _GEN_514 = !_T_893 ? sectored_entries_4_valid_2
			: _T_915 ? sectored_entries_4_valid_2 
			: _T_932 ? sectored_entries_4_valid_2 
			: _T_1062 ? _GEN_174 
			: sectored_entries_4_valid_2;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_4_valid_2 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2846 & sectored_entries_4_data_2[0]) begin
				    sectored_entries_4_valid_2 <= 1'h0;
				end else begin
					if (_T_406 & (2'h0 == _T_477)) begin
						sectored_entries_4_valid_2 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1062) begin
							sectored_entries_4_valid_2 <= _GEN_174;
						end
					end
				end
			end else begin
				sectored_entries_4_valid_2 <= io_sfence_bits_rs2 & (!sectored_entries_4_data_2[12] ? 1'h0 : _GEN_514);
			end
		end else begin
			sectored_entries_4_valid_2 <= _GEN_514;
		end
	end
end

  wire _GEN_175 = _GEN_953 
		| (_T_995 ? 1'h0 : sectored_entries_4_valid_3);
  wire _GEN_515 = !_T_893 ? sectored_entries_4_valid_3
			: _T_915 ? sectored_entries_4_valid_3 
			: _T_932 ? sectored_entries_4_valid_3 
			: _T_1062 ? _GEN_175 
			: sectored_entries_4_valid_3;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_4_valid_3 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2846 & sectored_entries_4_data_3[0]) begin
				    sectored_entries_4_valid_3 <= 1'h0;
				end else begin
					if (_T_406 & (2'h0 == _T_477)) begin
						sectored_entries_4_valid_3 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1062) begin
							sectored_entries_4_valid_3 <= _GEN_175;
						end
					end
				end
			end else begin
				sectored_entries_4_valid_3 <= io_sfence_bits_rs2 & (!sectored_entries_4_data_3[12] ? 1'h0 : _GEN_515);
			end
		end else begin
			sectored_entries_4_valid_3 <= _GEN_515;
		end
	end
end
// Passed
  wire _T_1079 = _T_993 == 3'h5;
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & !(_T_932) & _T_1079) begin
		sectored_entries_5_tag <= r_refill_tag;
		if (2'h0 == r_refill_tag[1:0]) begin
			sectored_entries_5_data_0 <= _T_931;
		end
		if (2'h1 == r_refill_tag[1:0]) begin
			sectored_entries_5_data_1 <= _T_931;
		end
		if (2'h2 == r_refill_tag[1:0]) begin
			sectored_entries_5_data_2 <= _T_931;
		end
		if (2'h3 == r_refill_tag[1:0]) begin
			sectored_entries_5_data_3 <= _T_931;
		end
	end
end

  wire _T_2993 = _T_410[19:10] == 10'h0;
  wire _GEN_194 = _GEN_950 
		| (_T_995 ? 1'h0 : sectored_entries_5_valid_0);
  wire _GEN_522 = !_T_893 ? sectored_entries_5_valid_0
			: _T_915 ? sectored_entries_5_valid_0 
			: _T_932 ? sectored_entries_5_valid_0 
			: _T_1079 ? _GEN_194 
			: sectored_entries_5_valid_0;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_5_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2993 & sectored_entries_5_data_0[0]) begin
				    sectored_entries_5_valid_0 <= 1'h0;
				end else begin
					if (_T_412 & (2'h0 == _T_477)) begin
						sectored_entries_5_valid_0 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1079) begin
							sectored_entries_5_valid_0 <= _GEN_194;
						end
					end
				end
			end else begin
				sectored_entries_5_valid_0 <= io_sfence_bits_rs2 & (!sectored_entries_5_data_0[12] ? 1'h0 : _GEN_522);
			end
		end else begin
			sectored_entries_5_valid_0 <= _GEN_522;
		end
	end
end

  wire _GEN_195 = _GEN_951 
		| (_T_995 ? 1'h0 : sectored_entries_5_valid_1);
  wire _GEN_523 = !_T_893 ? sectored_entries_5_valid_1
			: _T_915 ? sectored_entries_5_valid_1 
			: _T_932 ? sectored_entries_5_valid_1 
			: _T_1079 ? _GEN_195 
			: sectored_entries_5_valid_1;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_5_valid_1 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2993 & sectored_entries_5_data_1[0]) begin
				    sectored_entries_5_valid_1 <= 1'h0;
				end else begin
					if (_T_412 & (2'h0 == _T_477)) begin
						sectored_entries_5_valid_1 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1079) begin
							sectored_entries_5_valid_1 <= _GEN_195;
						end
					end
				end
			end else begin
				sectored_entries_5_valid_1 <= io_sfence_bits_rs2 & (!sectored_entries_5_data_1[12] ? 1'h0 : _GEN_523);
			end
		end else begin
			sectored_entries_5_valid_1 <= _GEN_523;
		end
	end
end

  wire _GEN_196 = _GEN_952 
		| (_T_995 ? 1'h0 : sectored_entries_5_valid_2);
  wire _GEN_524 = !_T_893 ? sectored_entries_5_valid_2
			: _T_915 ? sectored_entries_5_valid_2 
			: _T_932 ? sectored_entries_5_valid_2 
			: _T_1079 ? _GEN_196 
			: sectored_entries_5_valid_2;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_5_valid_2 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2993 & sectored_entries_5_data_2[0]) begin
				    sectored_entries_5_valid_2 <= 1'h0;
				end else begin
					if (_T_412 & (2'h0 == _T_477)) begin
						sectored_entries_5_valid_2 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1079) begin
							sectored_entries_5_valid_2 <= _GEN_196;
						end
					end
				end
			end else begin
				sectored_entries_5_valid_2 <= io_sfence_bits_rs2 & (!sectored_entries_5_data_2[12] ? 1'h0 : _GEN_524);
			end
		end else begin
			sectored_entries_5_valid_2 <= _GEN_524;
		end
	end
end

  wire _GEN_197 = _GEN_953 
		| (_T_995 ? 1'h0 : sectored_entries_5_valid_3);
  wire _GEN_525 = !_T_893 ? sectored_entries_5_valid_3
			: _T_915 ? sectored_entries_5_valid_3 
			: _T_932 ? sectored_entries_5_valid_3 
			: _T_1079 ? _GEN_197 
			: sectored_entries_5_valid_3;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_5_valid_3 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_2993 & sectored_entries_5_data_3[0]) begin
				    sectored_entries_5_valid_3 <= 1'h0;
				end else begin
					if (_T_412 & (2'h0 == _T_477)) begin
						sectored_entries_5_valid_3 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1079) begin
							sectored_entries_5_valid_3 <= _GEN_197;
						end
					end
				end
			end else begin
				sectored_entries_5_valid_3 <= io_sfence_bits_rs2 & (!sectored_entries_5_data_3[12] ? 1'h0 : _GEN_525);
			end
		end else begin
			sectored_entries_5_valid_3 <= _GEN_525;
		end
	end
end

  wire _T_1096 = _T_993 == 3'h6;
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & !(_T_932) & _T_1096) begin
		sectored_entries_6_tag <= r_refill_tag;
		if (2'h0 == r_refill_tag[1:0]) begin
			sectored_entries_6_data_0 <= _T_931;
		end
		if (2'h1 == r_refill_tag[1:0]) begin
			sectored_entries_6_data_1 <= _T_931;
		end
		if (2'h2 == r_refill_tag[1:0]) begin
			sectored_entries_6_data_2 <= _T_931;
		end
		if (2'h3 == r_refill_tag[1:0]) begin
			sectored_entries_6_data_3 <= _T_931;
		end
	end
end

  wire _T_3140 = _T_416[19:10] == 10'h0;
  wire _GEN_216 = _GEN_950 
		| (_T_995 ? 1'h0 : sectored_entries_6_valid_0);
  wire _GEN_532 = !_T_893 ? sectored_entries_6_valid_0
			: _T_915 ? sectored_entries_6_valid_0 
			: _T_932 ? sectored_entries_6_valid_0 
			: _T_1096 ? _GEN_216 
			: sectored_entries_6_valid_0;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_6_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_3140 & sectored_entries_6_data_0[0]) begin
				    sectored_entries_6_valid_0 <= 1'h0;
				end else begin
					if (_T_418 & (2'h0 == _T_477)) begin
						sectored_entries_6_valid_0 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1096) begin
							sectored_entries_6_valid_0 <= _GEN_216;
						end
					end
				end
			end else begin
				sectored_entries_6_valid_0 <= io_sfence_bits_rs2 & (!sectored_entries_6_data_0[12] ? 1'h0 : _GEN_532);
			end
		end else begin
			sectored_entries_6_valid_0 <= _GEN_532;
		end
	end
end

  wire _GEN_217 = _GEN_951 
		| (_T_995 ? 1'h0 : sectored_entries_6_valid_1);
  wire _GEN_533 = !_T_893 ? sectored_entries_6_valid_1
			: _T_915 ? sectored_entries_6_valid_1 
			: _T_932 ? sectored_entries_6_valid_1 
			: _T_1096 ? _GEN_217 
			: sectored_entries_6_valid_1;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_6_valid_1 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_3140 & sectored_entries_6_data_1[0]) begin
				    sectored_entries_6_valid_1 <= 1'h0;
				end else begin
					if (_T_418 & (2'h0 == _T_477)) begin
						sectored_entries_6_valid_1 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1096) begin
							sectored_entries_6_valid_1 <= _GEN_217;
						end
					end
				end
			end else begin
				sectored_entries_6_valid_1 <= io_sfence_bits_rs2 & (!sectored_entries_6_data_1[12] ? 1'h0 : _GEN_533);
			end
		end else begin
			sectored_entries_6_valid_1 <= _GEN_533;
		end
	end
end

  wire _GEN_218 = _GEN_952 
		| (_T_995 ? 1'h0 : sectored_entries_6_valid_2);
  wire _GEN_534 = !_T_893 ? sectored_entries_6_valid_2
			: _T_915 ? sectored_entries_6_valid_2 
			: _T_932 ? sectored_entries_6_valid_2 
			: _T_1096 ? _GEN_218 
			: sectored_entries_6_valid_2;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_6_valid_2 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_3140 & sectored_entries_6_data_2[0]) begin
				    sectored_entries_6_valid_2 <= 1'h0;
				end else begin
					if (_T_418 & (2'h0 == _T_477)) begin
						sectored_entries_6_valid_2 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1096) begin
							sectored_entries_6_valid_2 <= _GEN_218;
						end
					end
				end
			end else begin
				sectored_entries_6_valid_2 <= io_sfence_bits_rs2 & (!sectored_entries_6_data_2[12] ? 1'h0 : _GEN_534);
			end
		end else begin
			sectored_entries_6_valid_2 <= _GEN_534;
		end
	end
end

  wire _GEN_219 = _GEN_953 
		| (_T_995 ? 1'h0 : sectored_entries_6_valid_3);
  wire _GEN_535 = !_T_893 ? sectored_entries_6_valid_3
			: _T_915 ? sectored_entries_6_valid_3 
			: _T_932 ? sectored_entries_6_valid_3 
			: _T_1096 ? _GEN_219 
			: sectored_entries_6_valid_3;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_6_valid_3 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_3140 & sectored_entries_6_data_3[0]) begin
				    sectored_entries_6_valid_3 <= 1'h0;
				end else begin
					if (_T_418 & (2'h0 == _T_477)) begin
						sectored_entries_6_valid_3 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1096) begin
							sectored_entries_6_valid_3 <= _GEN_219;
						end
					end
				end
			end else begin
				sectored_entries_6_valid_3 <= io_sfence_bits_rs2 & (!sectored_entries_6_data_3[12] ? 1'h0 : _GEN_535);
			end
		end else begin
			sectored_entries_6_valid_3 <= _GEN_535;
		end
	end
end

  wire _T_1113 = _T_993 == 3'h7;
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & !(_T_932) & _T_1113) begin
		sectored_entries_7_tag <= r_refill_tag;
		if (2'h0 == r_refill_tag[1:0]) begin
			sectored_entries_7_data_0 <= _T_931;
		end
		if (2'h1 == r_refill_tag[1:0]) begin
			sectored_entries_7_data_1 <= _T_931;
		end
		if (2'h2 == r_refill_tag[1:0]) begin
			sectored_entries_7_data_2 <= _T_931;
		end
		if (2'h3 == r_refill_tag[1:0]) begin
			sectored_entries_7_data_3 <= _T_931;
		end
	end
end

  wire _T_3287 = _T_422[19:10] == 10'h0;
  wire _GEN_238 = _GEN_950 
		| (_T_995 ? 1'h0 : sectored_entries_7_valid_0);
  wire _GEN_542 = !_T_893 ? sectored_entries_7_valid_0
			: _T_915 ? sectored_entries_7_valid_0 
			: _T_932 ? sectored_entries_7_valid_0 
			: _T_1113 ? _GEN_238 
			: sectored_entries_7_valid_0;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_7_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_3287 & sectored_entries_7_data_0[0]) begin
				    sectored_entries_7_valid_0 <= 1'h0;
				end else begin
					if (_T_424 & (2'h0 == _T_477)) begin
						sectored_entries_7_valid_0 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1113) begin
							sectored_entries_7_valid_0 <= _GEN_238;
						end
					end
				end
			end else begin
				sectored_entries_7_valid_0 <= io_sfence_bits_rs2 & (!sectored_entries_7_data_0[12] ? 1'h0 : _GEN_542);
			end
		end else begin
			sectored_entries_7_valid_0 <= _GEN_542;
		end
	end
end

  wire _GEN_239 = _GEN_951 
		| (_T_995 ? 1'h0 : sectored_entries_7_valid_1);
  wire _GEN_543 = !_T_893 ? sectored_entries_7_valid_1
			: _T_915 ? sectored_entries_7_valid_1 
			: _T_932 ? sectored_entries_7_valid_1 
			: _T_1113 ? _GEN_239 
			: sectored_entries_7_valid_1;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_7_valid_1 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_3287 & sectored_entries_7_data_1[0]) begin
				    sectored_entries_7_valid_1 <= 1'h0;
				end else begin
					if (_T_424 & (2'h0 == _T_477)) begin
						sectored_entries_7_valid_1 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1113) begin
							sectored_entries_7_valid_1 <= _GEN_239;
						end
					end
				end
			end else begin
				sectored_entries_7_valid_1 <= io_sfence_bits_rs2 & (!sectored_entries_7_data_1[12] ? 1'h0 : _GEN_543);
			end
		end else begin
			sectored_entries_7_valid_1 <= _GEN_543;
		end
	end
end

  wire _GEN_240 = _GEN_952 
		| (_T_995 ? 1'h0 : sectored_entries_7_valid_2);
  wire _GEN_544 = !_T_893 ? sectored_entries_7_valid_2
			: _T_915 ? sectored_entries_7_valid_2 
			: _T_932 ? sectored_entries_7_valid_2 
			: _T_1113 ? _GEN_240 
			: sectored_entries_7_valid_2;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_7_valid_2 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_3287 & sectored_entries_7_data_2[0]) begin
				    sectored_entries_7_valid_2 <= 1'h0;
				end else begin
					if (_T_424 & (2'h0 == _T_477)) begin
						sectored_entries_7_valid_2 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1113) begin
							sectored_entries_7_valid_2 <= _GEN_240;
						end
					end
				end
			end else begin
				sectored_entries_7_valid_2 <= io_sfence_bits_rs2 & (!sectored_entries_7_data_2[12] ? 1'h0 : _GEN_544);
			end
		end else begin
			sectored_entries_7_valid_2 <= _GEN_544;
		end
	end
end

  wire _GEN_241 = _GEN_953 
		| (_T_995 ? 1'h0 : sectored_entries_7_valid_3);
  wire _GEN_545 = !_T_893 ? sectored_entries_7_valid_3
			: _T_915 ? sectored_entries_7_valid_3 
			: _T_932 ? sectored_entries_7_valid_3 
			: _T_1113 ? _GEN_241 
			: sectored_entries_7_valid_3;
always @(posedge clock) begin
	if (_T_3589) begin
		sectored_entries_7_valid_3 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_3287 & sectored_entries_7_data_3[0]) begin
				    sectored_entries_7_valid_3 <= 1'h0;
				end else begin
					if (_T_424 & (2'h0 == _T_477)) begin
						sectored_entries_7_valid_3 <= 1'h0;
					end else begin
						if (_T_893 & !(_T_915) & !(_T_932) & _T_1113) begin
							sectored_entries_7_valid_3 <= _GEN_241;
						end
					end
				end
			end else begin
				sectored_entries_7_valid_3 <= io_sfence_bits_rs2 & (!sectored_entries_7_data_3[12] ? 1'h0 : _GEN_545);
			end
		end else begin
			sectored_entries_7_valid_3 <= _GEN_545;
		end
	end
end
// Passed
  wire _T_933 = r_superpage_repl_addr == 2'h0;
  wire _T_948 = r_superpage_repl_addr == 2'h1;
  wire _T_963 = r_superpage_repl_addr == 2'h2;
  wire _T_978 = r_superpage_repl_addr == 2'h3;
  wire _GEN_66 = _T_933 | superpage_entries_0_valid_0;
  wire _GEN_70 = _T_948 | superpage_entries_1_valid_0;
  wire _GEN_74 = _T_963 | superpage_entries_2_valid_0;
  wire _GEN_78 = _T_978 | superpage_entries_3_valid_0;
  wire _GEN_858 = io_sfence_bits_rs2 & 
		(!superpage_entries_0_data_0[12] ? 1'h0 
		: !_T_893 ? superpage_entries_0_valid_0 
		: _T_915 ? superpage_entries_0_valid_0 
		: _T_932 ? _GEN_66 
		: superpage_entries_0_valid_0
		);
  wire _GEN_862 = io_sfence_bits_rs2 & 
		(!superpage_entries_1_data_0[12] ? 1'h0 
		: !_T_893 ? superpage_entries_1_valid_0 
		: _T_915 ? superpage_entries_1_valid_0 
		: _T_932 ? _GEN_70 
		: superpage_entries_1_valid_0
		);
  wire _GEN_866 = io_sfence_bits_rs2 & 
		(!superpage_entries_2_data_0[12] ? 1'h0 
		: !_T_893 ? superpage_entries_2_valid_0
		: _T_915 ? superpage_entries_2_valid_0 
		: _T_932 ? _GEN_74 
		: superpage_entries_2_valid_0
		);
  wire _GEN_870 = io_sfence_bits_rs2 & 
		(!superpage_entries_3_data_0[12] ? 1'h0 
		: !_T_893 ? superpage_entries_3_valid_0
		: _T_915 ? superpage_entries_3_valid_0 
		: _T_932 ? _GEN_78 
		: superpage_entries_3_valid_0
		); 
always @(posedge clock) begin
	if (_T_893 & !(_T_915) & _T_932) begin
		if (_T_933) begin
			superpage_entries_0_tag <= r_refill_tag;
			superpage_entries_0_data_0 <= _T_931;
		end
		if (_T_948) begin
			superpage_entries_1_tag <= r_refill_tag;
			superpage_entries_1_data_0 <= _T_931;
		end
		if (_T_963) begin
			superpage_entries_2_tag <= r_refill_tag;
			superpage_entries_2_data_0 <= _T_931;
		end
		if (_T_978) begin
			superpage_entries_3_tag <= r_refill_tag;
			superpage_entries_3_data_0 <= _T_931;
		end
	end
	if (_T_3589) begin
		superpage_entries_0_valid_0 <= 1'h0;
		superpage_entries_1_valid_0 <= 1'h0;
		superpage_entries_2_valid_0 <= 1'h0;
		superpage_entries_3_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (superpage_hits_0) begin
					superpage_entries_0_valid_0 <= 1'h0;
				end else begin
					if (_T_893 & !(_T_915) & _T_932) begin
						superpage_entries_0_valid_0 <= _GEN_66;
					end
				end
				if (superpage_hits_1) begin
					superpage_entries_1_valid_0 <= 1'h0;
				end else begin
					if (_T_893 & !(_T_915) & _T_932) begin
				        	superpage_entries_1_valid_0 <= _GEN_70;
					end
				end
				if (superpage_hits_2) begin
					superpage_entries_2_valid_0 <= 1'h0;
				end else begin
					if (_T_893 & !(_T_915) & _T_932) begin
				        	superpage_entries_2_valid_0 <= _GEN_74;
					end
				end
				if (superpage_hits_3) begin
					superpage_entries_3_valid_0 <= 1'h0;
				end else begin
					if (_T_893 & !(_T_915) & _T_932) begin
				        	superpage_entries_3_valid_0 <= _GEN_78;
					end
				end
			end else begin
				superpage_entries_0_valid_0 <= _GEN_858;
				superpage_entries_1_valid_0 <= _GEN_862;
				superpage_entries_2_valid_0 <= _GEN_866;
				superpage_entries_3_valid_0 <= _GEN_870;
			end
		end else begin
			if (_T_893 & !(_T_915) & _T_932) begin
				superpage_entries_0_valid_0 <= _GEN_66;
				superpage_entries_1_valid_0 <= _GEN_70;
				superpage_entries_2_valid_0 <= _GEN_74;
				superpage_entries_3_valid_0 <= _GEN_78;
			end
		end
	end
end

  wire _GEN_354 = _T_915 | special_entry_valid_0;
  wire _GEN_874 = io_sfence_bits_rs2 & 
		(!special_entry_data_0[12] ? 1'h0 
		: !_T_893 ? special_entry_valid_0
		: _GEN_354
		);
always @(posedge clock) begin
	if (_T_893 & _T_915) begin
		special_entry_level <= io_ptw_resp_bits_level;
		special_entry_tag <= r_refill_tag;
		special_entry_data_0 <= _T_931;
	end
	if (_T_3589) begin
		special_entry_valid_0 <= 1'h0;
	end else begin
		if (io_sfence_valid) begin
			if (io_sfence_bits_rs1) begin
				if (_T_586) begin
					special_entry_valid_0 <= 1'h0;
				end else begin
					if (_T_893) begin
						special_entry_valid_0 <= _GEN_354;
					end
				end
			end else begin
				special_entry_valid_0 <= _GEN_874;
			end
		end else begin
			if (_T_893) begin
				special_entry_valid_0 <= _GEN_354;
			end
		end
	end
end

  wire _T_2114 = io_req_ready & io_req_valid & tlb_miss;
always @(posedge clock) begin
	if (reset) begin
		state <= 2'h0;
	end else begin
		if (io_ptw_resp_valid) begin
			state <= 2'h0;
		end else begin
			if ((state == 2'h2) & io_sfence_valid) begin
				state <= 2'h3;
			end else begin
				if (_T_4) begin
					if (io_ptw_req_ready) begin
						if (io_sfence_valid) begin
							state <= 2'h3;
						end else begin
							state <= 2'h2;
						end
					end else begin
						if (io_sfence_valid) begin
							state <= 2'h0;
						end else begin
							if (_T_2114) begin
								state <= 2'h1;
							end
						end
					end
				end else begin
					if (_T_2114) begin
						state <= 2'h1;
					end
				end
			end
		end
	end
end

  wire [3:0] _T_2126 = {_T_1905, 1'h0} >> {1'h1,_T_1905[0]};
always @(posedge clock) begin
	if (_T_2114) begin
		r_refill_tag <= vpn;
	end
	if (_T_2114) begin
		if ({superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0} == 4'hf) begin
			r_superpage_repl_addr <= {_T_1905[0],_T_2126[0]};
		end else begin
			if (!superpage_entries_0_valid_0) begin
				r_superpage_repl_addr <= 2'h0;
			end else begin
				if (!superpage_entries_1_valid_0) begin
					r_superpage_repl_addr <= 2'h1;
				end else begin
					if (!superpage_entries_2_valid_0) begin
						r_superpage_repl_addr <= 2'h2;
					end else begin
						r_superpage_repl_addr <= 2'h3;
					end
				end
			end
		end
	end
end

  wire _T_1913 = sector_hits_0 
		| sector_hits_1 
		| sector_hits_2 
		| sector_hits_3 
		| sector_hits_4 
		| sector_hits_5 
		| sector_hits_6 
		| sector_hits_7;
  wire [7:0] _T_1920 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0};
  wire _T_1923 = _T_1920[7:4] != 4'h0;
  wire [3:0] _T_1924 = _T_1920[7:4] | _T_1920[3:0];
  wire _T_1927 = _T_1924[3:2] != 2'h0;
  wire [1:0] _T_1928 = _T_1924[3:2] | _T_1924[1:0];
  wire [2:0] _T_1931 = {_T_1923,_T_1927,_T_1928[1]};
  wire [7:0] _T_1932 = {_T_1904, 1'h0};
  wire [7:0] _T_2148 = {{1'd0}, _T_1932[7:1]};
  wire [7:0] _T_2155 = _T_1932 >> {1'h1,_T_2148[0]};
  wire [7:0] _T_2162 = _T_1932 >> {1'h1,_T_2148[0],_T_2155[0]};
  wire [3:0] _T_2165 = {1'h1,_T_2148[0],_T_2155[0],_T_2162[0]}; 
always @(posedge clock) begin
	if (_T_2114) begin
		if ({_T_421,_T_415,_T_409,_T_403,_T_397,_T_391,_T_385,_T_379} == 8'hff) begin
			r_sectored_repl_addr <= _T_2165[2:0];
		end else if (!_T_379) begin
			r_sectored_repl_addr <= 3'h0;
		end else if (!_T_385) begin
			r_sectored_repl_addr <= 3'h1;
		end else if (!_T_391) begin
			r_sectored_repl_addr <= 3'h2;
		end else if (!_T_397) begin
			r_sectored_repl_addr <= 3'h3;
		end else if (!_T_403) begin
			r_sectored_repl_addr <= 3'h4;
		end else if (!_T_409) begin
			r_sectored_repl_addr <= 3'h5;
		end else if (!_T_415) begin
			r_sectored_repl_addr <= 3'h6;
		end else begin
			r_sectored_repl_addr <= 3'h7;
		end
	end
	if (_T_2114) begin
		r_sectored_hit_addr <= _T_1931;
	end
	if (_T_2114) begin
		r_sectored_hit <= _T_1913;
	end
end

  wire [7:0] _T_1940 = !_T_1931[2] ? (_T_1932 | 8'h2) : ~ ((~ _T_1932) | 8'h2);
  wire [3:0] _T_1944 = 4'h1 << {1'h1,_T_1931[2]};
  wire [7:0] _T_1949 = !_T_1931[1] ? (_T_1940 | {{4'd0}, _T_1944}) : (~ ((~ _T_1940) | {{4'd0}, _T_1944}));
  wire [7:0] _T_1953 = 8'h1 << {1'h1,_T_1931[2],_T_1931[1]};
  wire [7:0] _T_1958 = !_T_1931[0] ? (_T_1949 | _T_1953) : (~ ((~ _T_1949) | _T_1953));
  wire [3:0] _T_1966 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0};
  wire _T_1969 = _T_1966[3:2] != 2'h0;
  wire [1:0] _T_1970 = _T_1966[3:2] | _T_1966[1:0];
  wire [1:0] _T_1972 = {_T_1969,_T_1970[1]};
  wire [3:0] _T_1981 = !_T_1972[1] ? ({_T_1905, 1'h0} | 4'h2) : (~ ((~ {_T_1905, 1'h0}) | 4'h2));
  wire [3:0] _T_1985 = 4'h1 << {1'h1,_T_1972[1]};
  wire [3:0] _T_1990 = !_T_1972[0] ? (_T_1981 | _T_1985) : (~ ((~ _T_1981) | _T_1985));
always @(posedge clock) begin
	if (io_req_valid & vm_enabled) begin
		if (_T_1913) begin
			_T_1904 <= _T_1958[7:1];
		end
		if (superpage_hits_0 | superpage_hits_1 | superpage_hits_2 | superpage_hits_3) begin
			_T_1905 <= _T_1990[3:1];
		end
	end
end

  wire _T_2251 = (!io_sfence_bits_rs1 | (io_sfence_bits_addr[31:12] == vpn) | reset) == 1'h0;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & _T_2251) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:368 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & _T_2251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_72[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_73[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_75[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_76[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_78[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_79[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_81[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_82[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  special_entry_level = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  special_entry_tag = _RAND_85[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_86[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  state = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  r_refill_tag = _RAND_89[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_90[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_92[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_sectored_hit = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1904 = _RAND_94[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1905 = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end

`endif // MY_ASSIGNMENT

endmodule
`endif // __TLB

