`include "include_module.v"
`ifdef __TLB_1
module TLB_1( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129454.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129455.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129456.4]
  output        io_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_req_bits_vaddr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  output        io_resp_miss, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  output [31:0] io_resp_paddr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  output        io_resp_pf_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  output        io_resp_ae_inst, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  output        io_resp_cacheable, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_sfence_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_sfence_bits_rs1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_sfence_bits_rs2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_sfence_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  output        io_ptw_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  output        io_ptw_req_bits_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  output [19:0] io_ptw_req_bits_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_ae, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [53:0] io_ptw_resp_bits_pte_ppn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_pte_d, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_pte_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_pte_g, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_pte_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_pte_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_pte_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_pte_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_pte_v, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_level, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_resp_bits_homogeneous, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_ptbr_mode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_status_debug, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_status_prv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_0_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_pmp_0_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_0_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_0_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_0_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [29:0] io_ptw_pmp_0_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_ptw_pmp_0_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_1_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_pmp_1_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_1_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_1_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_1_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [29:0] io_ptw_pmp_1_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_ptw_pmp_1_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_2_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_pmp_2_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_2_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_2_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_2_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [29:0] io_ptw_pmp_2_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_ptw_pmp_2_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_3_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_pmp_3_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_3_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_3_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_3_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [29:0] io_ptw_pmp_3_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_ptw_pmp_3_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_4_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_pmp_4_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_4_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_4_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_4_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [29:0] io_ptw_pmp_4_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_ptw_pmp_4_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_5_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_pmp_5_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_5_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_5_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_5_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [29:0] io_ptw_pmp_5_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_ptw_pmp_5_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_6_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_pmp_6_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_6_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_6_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_6_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [29:0] io_ptw_pmp_6_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_ptw_pmp_6_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_7_cfg_l, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [1:0]  io_ptw_pmp_7_cfg_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_7_cfg_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_7_cfg_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_ptw_pmp_7_cfg_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [29:0] io_ptw_pmp_7_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input  [31:0] io_ptw_pmp_7_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
  input         io_kill // @[:freechips.rocketchip.system.DefaultRV32Config.fir@129457.4]
);
  wire [19:0] _2_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire [19:0] _2_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire  _2_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
  wire [1:0] pmp_io_prv; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [31:0] pmp_io_addr; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_r; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_w; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire  pmp_io_x; // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
  wire [19:0] _2_1_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire [19:0] _2_1_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire  _2_1_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
  wire [19:0] _2_2_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire [19:0] _2_2_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire  _2_2_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
  wire [19:0] _2_3_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire [19:0] _2_3_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire  _2_3_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
  wire [19:0] _2_4_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire [19:0] _2_4_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire  _2_4_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
  wire [19:0] _2_5_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire [19:0] _2_5_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire  _2_5_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
  wire [19:0] _2_6_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire [19:0] _2_6_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire  _2_6_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
  wire [19:0] _2_7_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire [19:0] _2_7_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire  _2_7_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
  wire [19:0] _2_8_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire [19:0] _2_8_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire  _2_8_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
  wire [19:0] _2_9_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire [19:0] _2_9_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire  _2_9_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
  wire [19:0] _2_10_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire [19:0] _2_10_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire  _2_10_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
  wire [19:0] _2_11_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire [19:0] _2_11_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire  _2_11_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
  wire [19:0] _2_12_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire [19:0] _2_12_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire  _2_12_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
  wire [19:0] _2_13_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire [19:0] _2_13_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire  _2_13_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
  wire [19:0] _2_14_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire [19:0] _2_14_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire  _2_14_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
  wire [19:0] _2_15_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire [19:0] _2_15_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire  _2_15_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
  wire [19:0] _2_16_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire [19:0] _2_16_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire  _2_16_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
  wire [19:0] _2_17_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire [19:0] _2_17_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire  _2_17_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
  wire [19:0] _2_18_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire [19:0] _2_18_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire  _2_18_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
  wire [19:0] _2_19_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire [19:0] _2_19_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire  _2_19_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
  wire [19:0] _2_20_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire [19:0] _2_20_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire  _2_20_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
  wire [19:0] _2_21_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire [19:0] _2_21_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire  _2_21_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
  wire [19:0] _2_22_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire [19:0] _2_22_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire  _2_22_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
  wire [19:0] _2_23_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire [19:0] _2_23_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire  _2_23_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
  wire [19:0] _2_24_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire [19:0] _2_24_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire  _2_24_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
  wire [19:0] _2_25_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire [19:0] _2_25_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire  _2_25_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
  wire [19:0] _2_26_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire [19:0] _2_26_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire  _2_26_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
  wire [19:0] _2_27_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire [19:0] _2_27_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire  _2_27_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
  wire [19:0] _2_28_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire [19:0] _2_28_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire  _2_28_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
  wire [19:0] _2_29_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire [19:0] _2_29_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire  _2_29_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
  wire [19:0] _2_30_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire [19:0] _2_30_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire  _2_30_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
  wire [19:0] _2_31_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire [19:0] _2_31_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire  _2_31_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
  wire [19:0] _2_32_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire [19:0] _2_32_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire  _2_32_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
  wire [19:0] _2_33_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire [19:0] _2_33_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire  _2_33_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
  wire [19:0] _2_34_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire [19:0] _2_34_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire  _2_34_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
  wire [19:0] _2_35_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire [19:0] _2_35_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire  _2_35_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
  wire [19:0] _2_36_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire [19:0] _2_36_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire  _2_36_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
  wire [19:0] _2_37_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire [19:0] _2_37_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire  _2_37_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
  wire [19:0] _2_38_io_x_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_x_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire [19:0] _2_38_io_y_ppn; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_u; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_ae; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_sw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_sx; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_sr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_pw; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_px; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_pr; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_pal; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_paa; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_eff; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  wire  _2_38_io_y_c; // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
  reg [19:0] sectored_entries_0_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_0;
  reg [33:0] sectored_entries_0_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_1;
  reg [33:0] sectored_entries_0_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_2;
  reg [33:0] sectored_entries_0_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_3;
  reg [33:0] sectored_entries_0_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_8;
  reg [19:0] sectored_entries_1_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_9;
  reg [33:0] sectored_entries_1_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_10;
  reg [33:0] sectored_entries_1_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_11;
  reg [33:0] sectored_entries_1_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_12;
  reg [33:0] sectored_entries_1_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_13;
  reg  sectored_entries_1_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_14;
  reg  sectored_entries_1_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_15;
  reg  sectored_entries_1_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_16;
  reg  sectored_entries_1_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_17;
  reg [19:0] sectored_entries_2_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_18;
  reg [33:0] sectored_entries_2_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_19;
  reg [33:0] sectored_entries_2_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_20;
  reg [33:0] sectored_entries_2_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_21;
  reg [33:0] sectored_entries_2_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_22;
  reg  sectored_entries_2_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_23;
  reg  sectored_entries_2_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_24;
  reg  sectored_entries_2_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_25;
  reg  sectored_entries_2_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_26;
  reg [19:0] sectored_entries_3_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_27;
  reg [33:0] sectored_entries_3_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_28;
  reg [33:0] sectored_entries_3_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_29;
  reg [33:0] sectored_entries_3_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_30;
  reg [33:0] sectored_entries_3_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_31;
  reg  sectored_entries_3_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_32;
  reg  sectored_entries_3_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_33;
  reg  sectored_entries_3_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_34;
  reg  sectored_entries_3_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_35;
  reg [19:0] sectored_entries_4_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_36;
  reg [33:0] sectored_entries_4_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_37;
  reg [33:0] sectored_entries_4_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_38;
  reg [33:0] sectored_entries_4_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_39;
  reg [33:0] sectored_entries_4_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_40;
  reg  sectored_entries_4_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_41;
  reg  sectored_entries_4_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_42;
  reg  sectored_entries_4_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_43;
  reg  sectored_entries_4_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_44;
  reg [19:0] sectored_entries_5_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_45;
  reg [33:0] sectored_entries_5_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_46;
  reg [33:0] sectored_entries_5_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_47;
  reg [33:0] sectored_entries_5_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_48;
  reg [33:0] sectored_entries_5_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_49;
  reg  sectored_entries_5_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_50;
  reg  sectored_entries_5_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_51;
  reg  sectored_entries_5_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_52;
  reg  sectored_entries_5_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_53;
  reg [19:0] sectored_entries_6_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_54;
  reg [33:0] sectored_entries_6_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_55;
  reg [33:0] sectored_entries_6_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_56;
  reg [33:0] sectored_entries_6_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_57;
  reg [33:0] sectored_entries_6_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_58;
  reg  sectored_entries_6_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_59;
  reg  sectored_entries_6_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_60;
  reg  sectored_entries_6_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_61;
  reg  sectored_entries_6_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_62;
  reg [19:0] sectored_entries_7_tag; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_63;
  reg [33:0] sectored_entries_7_data_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_64;
  reg [33:0] sectored_entries_7_data_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_65;
  reg [33:0] sectored_entries_7_data_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_66;
  reg [33:0] sectored_entries_7_data_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [63:0] _RAND_67;
  reg  sectored_entries_7_valid_0; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_68;
  reg  sectored_entries_7_valid_1; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_69;
  reg  sectored_entries_7_valid_2; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_70;
  reg  sectored_entries_7_valid_3; // @[TLB.scala 161:29:freechips.rocketchip.system.DefaultRV32Config.fir@129462.4]
  reg [31:0] _RAND_71;
  reg [19:0] superpage_entries_0_tag; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [31:0] _RAND_72;
  reg [33:0] superpage_entries_0_data_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [63:0] _RAND_73;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [31:0] _RAND_74;
  reg [19:0] superpage_entries_1_tag; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [31:0] _RAND_75;
  reg [33:0] superpage_entries_1_data_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [63:0] _RAND_76;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [31:0] _RAND_77;
  reg [19:0] superpage_entries_2_tag; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [31:0] _RAND_78;
  reg [33:0] superpage_entries_2_data_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [63:0] _RAND_79;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [31:0] _RAND_80;
  reg [19:0] superpage_entries_3_tag; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [31:0] _RAND_81;
  reg [33:0] superpage_entries_3_data_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [63:0] _RAND_82;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 162:30:freechips.rocketchip.system.DefaultRV32Config.fir@129463.4]
  reg [31:0] _RAND_83;
  reg  special_entry_level; // @[TLB.scala 163:56:freechips.rocketchip.system.DefaultRV32Config.fir@129464.4]
  reg [31:0] _RAND_84;
  reg [19:0] special_entry_tag; // @[TLB.scala 163:56:freechips.rocketchip.system.DefaultRV32Config.fir@129464.4]
  reg [31:0] _RAND_85;
  reg [33:0] special_entry_data_0; // @[TLB.scala 163:56:freechips.rocketchip.system.DefaultRV32Config.fir@129464.4]
  reg [63:0] _RAND_86;
  reg  special_entry_valid_0; // @[TLB.scala 163:56:freechips.rocketchip.system.DefaultRV32Config.fir@129464.4]
  reg [31:0] _RAND_87;
  reg [1:0] state; // @[TLB.scala 168:18:freechips.rocketchip.system.DefaultRV32Config.fir@129465.4]
  reg [31:0] _RAND_88;
  reg [19:0] r_refill_tag; // @[TLB.scala 169:25:freechips.rocketchip.system.DefaultRV32Config.fir@129466.4]
  reg [31:0] _RAND_89;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 170:34:freechips.rocketchip.system.DefaultRV32Config.fir@129467.4]
  reg [31:0] _RAND_90;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 171:33:freechips.rocketchip.system.DefaultRV32Config.fir@129468.4]
  reg [31:0] _RAND_91;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 172:32:freechips.rocketchip.system.DefaultRV32Config.fir@129469.4]
  reg [31:0] _RAND_92;
  reg  r_sectored_hit; // @[TLB.scala 173:27:freechips.rocketchip.system.DefaultRV32Config.fir@129470.4]
  reg [31:0] _RAND_93;
  wire  priv_s; // @[TLB.scala 176:20:freechips.rocketchip.system.DefaultRV32Config.fir@129471.4]
  wire  priv_uses_vm; // @[TLB.scala 177:27:freechips.rocketchip.system.DefaultRV32Config.fir@129472.4]
  wire  vm_enabled; // @[TLB.scala 178:83:freechips.rocketchip.system.DefaultRV32Config.fir@129475.4]
  wire [19:0] vpn; // @[TLB.scala 181:30:freechips.rocketchip.system.DefaultRV32Config.fir@129478.4]
  wire [19:0] refill_ppn; // @[TLB.scala 182:44:freechips.rocketchip.system.DefaultRV32Config.fir@129479.4]
  wire  _T_4; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@129481.4]
  wire  _T_5; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@129482.4]
  wire  invalidate_refill; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129483.4]
  wire  _T_21; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@129514.4]
  wire [9:0] _T_24; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@129525.4]
  wire  _T_25; // @[TLB.scala 121:30:freechips.rocketchip.system.DefaultRV32Config.fir@129526.4]
  wire [19:0] _T_27; // @[TLB.scala 122:30:freechips.rocketchip.system.DefaultRV32Config.fir@129528.4]
  wire [19:0] _T_28; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@129529.4]
  wire [9:0] _T_29; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@129530.4]
  wire [19:0] _T_30; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@129531.4]
  wire [19:0] _T_31; // @[TLB.scala 186:123:freechips.rocketchip.system.DefaultRV32Config.fir@129532.4]
  wire [19:0] _T_32; // @[TLB.scala 186:20:freechips.rocketchip.system.DefaultRV32Config.fir@129533.4]
  wire [19:0] mpu_ppn; // @[TLB.scala 185:20:freechips.rocketchip.system.DefaultRV32Config.fir@129534.4]
  wire [11:0] _T_33; // @[TLB.scala 187:52:freechips.rocketchip.system.DefaultRV32Config.fir@129535.4]
  wire [31:0] mpu_physaddr; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@129536.4]
  wire [2:0] _T_36; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@129539.4]
  wire [2:0] mpu_priv; // @[TLB.scala 188:27:freechips.rocketchip.system.DefaultRV32Config.fir@129540.4]
  wire [31:0] _T_37; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129556.4]
  wire [32:0] _T_38; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129557.4]
  wire [32:0] _T_39; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129558.4]
  wire [32:0] _T_40; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129559.4]
  wire  _T_41; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129560.4]
  wire [31:0] _T_42; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129561.4]
  wire [32:0] _T_43; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129562.4]
  wire [32:0] _T_44; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129563.4]
  wire [32:0] _T_45; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129564.4]
  wire  _T_46; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129565.4]
  wire [31:0] _T_47; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129566.4]
  wire [32:0] _T_48; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129567.4]
  wire [32:0] _T_49; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129568.4]
  wire [32:0] _T_50; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129569.4]
  wire  _T_51; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129570.4]
  wire [32:0] _T_53; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129572.4]
  wire [32:0] _T_54; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129573.4]
  wire [32:0] _T_55; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129574.4]
  wire  _T_56; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129575.4]
  wire [31:0] _T_57; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129576.4]
  wire [32:0] _T_58; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129577.4]
  wire [32:0] _T_59; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129578.4]
  wire [32:0] _T_60; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129579.4]
  wire  _T_61; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129580.4]
  wire [31:0] _T_62; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129581.4]
  wire [32:0] _T_63; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129582.4]
  wire [32:0] _T_64; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129583.4]
  wire [32:0] _T_65; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129584.4]
  wire  _T_66; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129585.4]
  wire [31:0] _T_67; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129586.4]
  wire [32:0] _T_68; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129587.4]
  wire [32:0] _T_69; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129588.4]
  wire [32:0] _T_70; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129589.4]
  wire  _T_71; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129590.4]
  wire  _T_73; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129600.4]
  wire  _T_74; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129601.4]
  wire  _T_75; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129602.4]
  wire  _T_76; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129603.4]
  wire  _T_77; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129604.4]
  wire  legal_address; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129605.4]
  wire [32:0] _T_85; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129613.4]
  wire [32:0] _T_86; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129614.4]
  wire  _T_87; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129615.4]
  wire  cacheable; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129621.4]
  wire [31:0] _T_142; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129673.4]
  wire [32:0] _T_143; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129674.4]
  wire [32:0] _T_144; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129675.4]
  wire [32:0] _T_145; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129676.4]
  wire  _T_146; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129677.4]
  wire [32:0] _T_163; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129694.4]
  wire [32:0] _T_164; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129695.4]
  wire  _T_165; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129696.4]
  wire  _T_172; // @[TLBPermissions.scala 82:66:freechips.rocketchip.system.DefaultRV32Config.fir@129703.4]
  wire  _T_185; // @[TLB.scala 199:39:freechips.rocketchip.system.DefaultRV32Config.fir@129716.4]
  wire  deny_access_to_debug; // @[TLB.scala 199:48:freechips.rocketchip.system.DefaultRV32Config.fir@129722.4]
  wire  _T_197; // @[TLB.scala 200:44:freechips.rocketchip.system.DefaultRV32Config.fir@129729.4]
  wire  _T_198; // @[TLB.scala 200:41:freechips.rocketchip.system.DefaultRV32Config.fir@129730.4]
  wire  prot_r; // @[TLB.scala 200:66:freechips.rocketchip.system.DefaultRV32Config.fir@129731.4]
  wire [32:0] _T_211; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129744.4]
  wire [32:0] _T_212; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129745.4]
  wire  _T_213; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129746.4]
  wire [31:0] _T_214; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129747.4]
  wire [32:0] _T_215; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129748.4]
  wire [32:0] _T_216; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129749.4]
  wire [32:0] _T_217; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129750.4]
  wire  _T_218; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129751.4]
  wire  _T_220; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129753.4]
  wire  _T_221; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129754.4]
  wire  _T_231; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129765.4]
  wire  _T_233; // @[TLB.scala 201:45:freechips.rocketchip.system.DefaultRV32Config.fir@129767.4]
  wire  prot_w; // @[TLB.scala 201:70:freechips.rocketchip.system.DefaultRV32Config.fir@129768.4]
  wire  prot_al; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129802.4]
  wire [32:0] _T_300; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129839.4]
  wire [32:0] _T_301; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129840.4]
  wire  _T_302; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129841.4]
  wire  _T_313; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129852.4]
  wire  _T_314; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129853.4]
  wire  _T_330; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129870.4]
  wire  _T_332; // @[TLB.scala 204:40:freechips.rocketchip.system.DefaultRV32Config.fir@129872.4]
  wire  prot_x; // @[TLB.scala 204:65:freechips.rocketchip.system.DefaultRV32Config.fir@129873.4]
  wire [32:0] _T_357; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129898.4]
  wire [32:0] _T_358; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129899.4]
  wire  _T_359; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129900.4]
  wire [32:0] _T_362; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129903.4]
  wire [32:0] _T_363; // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129904.4]
  wire  _T_364; // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129905.4]
  wire  _T_370; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129911.4]
  wire  _T_371; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129912.4]
  wire  _T_372; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129913.4]
  wire  prot_eff; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129919.4]
  wire  _T_377; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129920.4]
  wire  _T_378; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129921.4]
  wire  _T_379; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129922.4]
  wire [19:0] _T_380; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129923.4]
  wire [17:0] _T_381; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129924.4]
  wire  _T_382; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129925.4]
  wire  sector_hits_0; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129926.4]
  wire  _T_383; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129927.4]
  wire  _T_384; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129928.4]
  wire  _T_385; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129929.4]
  wire [19:0] _T_386; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129930.4]
  wire [17:0] _T_387; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129931.4]
  wire  _T_388; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129932.4]
  wire  sector_hits_1; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129933.4]
  wire  _T_389; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129934.4]
  wire  _T_390; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129935.4]
  wire  _T_391; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129936.4]
  wire [19:0] _T_392; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129937.4]
  wire [17:0] _T_393; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129938.4]
  wire  _T_394; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129939.4]
  wire  sector_hits_2; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129940.4]
  wire  _T_395; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129941.4]
  wire  _T_396; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129942.4]
  wire  _T_397; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129943.4]
  wire [19:0] _T_398; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129944.4]
  wire [17:0] _T_399; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129945.4]
  wire  _T_400; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129946.4]
  wire  sector_hits_3; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129947.4]
  wire  _T_401; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129948.4]
  wire  _T_402; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129949.4]
  wire  _T_403; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129950.4]
  wire [19:0] _T_404; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129951.4]
  wire [17:0] _T_405; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129952.4]
  wire  _T_406; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129953.4]
  wire  sector_hits_4; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129954.4]
  wire  _T_407; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129955.4]
  wire  _T_408; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129956.4]
  wire  _T_409; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129957.4]
  wire [19:0] _T_410; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129958.4]
  wire [17:0] _T_411; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129959.4]
  wire  _T_412; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129960.4]
  wire  sector_hits_5; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129961.4]
  wire  _T_413; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129962.4]
  wire  _T_414; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129963.4]
  wire  _T_415; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129964.4]
  wire [19:0] _T_416; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129965.4]
  wire [17:0] _T_417; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129966.4]
  wire  _T_418; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129967.4]
  wire  sector_hits_6; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129968.4]
  wire  _T_419; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129969.4]
  wire  _T_420; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129970.4]
  wire  _T_421; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129971.4]
  wire [19:0] _T_422; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129972.4]
  wire [17:0] _T_423; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129973.4]
  wire  _T_424; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129974.4]
  wire  sector_hits_7; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129975.4]
  wire [9:0] _T_427; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@129978.4]
  wire [9:0] _T_428; // @[TLB.scala 108:86:freechips.rocketchip.system.DefaultRV32Config.fir@129979.4]
  wire  _T_429; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@129980.4]
  wire  superpage_hits_0; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@129982.4]
  wire [9:0] _T_435; // @[TLB.scala 108:86:freechips.rocketchip.system.DefaultRV32Config.fir@129986.4]
  wire [9:0] _T_440; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@129992.4]
  wire  _T_442; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@129994.4]
  wire  superpage_hits_1; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@129996.4]
  wire [9:0] _T_453; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@130006.4]
  wire  _T_455; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@130008.4]
  wire  superpage_hits_2; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@130010.4]
  wire [9:0] _T_466; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@130020.4]
  wire  _T_468; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@130022.4]
  wire  superpage_hits_3; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@130024.4]
  wire [1:0] _T_477; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@130032.4]
  wire  _GEN_1; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130036.4]
  wire  _GEN_2; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130036.4]
  wire  _GEN_3; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130036.4]
  wire  _T_481; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130036.4]
  wire  hitsVec_0; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130037.4]
  wire  _GEN_5; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130042.4]
  wire  _GEN_6; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130042.4]
  wire  _GEN_7; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130042.4]
  wire  _T_486; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130042.4]
  wire  hitsVec_1; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130043.4]
  wire  _GEN_9; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130048.4]
  wire  _GEN_10; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130048.4]
  wire  _GEN_11; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130048.4]
  wire  _T_491; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130048.4]
  wire  hitsVec_2; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130049.4]
  wire  _GEN_13; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130054.4]
  wire  _GEN_14; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130054.4]
  wire  _GEN_15; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130054.4]
  wire  _T_496; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130054.4]
  wire  hitsVec_3; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130055.4]
  wire  _GEN_17; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130060.4]
  wire  _GEN_18; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130060.4]
  wire  _GEN_19; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130060.4]
  wire  _T_501; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130060.4]
  wire  hitsVec_4; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130061.4]
  wire  _GEN_21; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130066.4]
  wire  _GEN_22; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130066.4]
  wire  _GEN_23; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130066.4]
  wire  _T_506; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130066.4]
  wire  hitsVec_5; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130067.4]
  wire  _GEN_25; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130072.4]
  wire  _GEN_26; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130072.4]
  wire  _GEN_27; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130072.4]
  wire  _T_511; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130072.4]
  wire  hitsVec_6; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130073.4]
  wire  _GEN_29; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130078.4]
  wire  _GEN_30; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130078.4]
  wire  _GEN_31; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130078.4]
  wire  _T_516; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130078.4]
  wire  hitsVec_7; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130079.4]
  wire  hitsVec_8; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130094.4]
  wire  hitsVec_9; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130109.4]
  wire  hitsVec_10; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130124.4]
  wire  hitsVec_11; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130139.4]
  wire [9:0] _T_575; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@130142.4]
  wire  _T_577; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@130144.4]
  wire  _T_579; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@130146.4]
  wire [9:0] _T_582; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@130149.4]
  wire  _T_584; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@130151.4]
  wire  _T_585; // @[TLB.scala 108:42:freechips.rocketchip.system.DefaultRV32Config.fir@130152.4]
  wire  _T_586; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@130153.4]
  wire  hitsVec_12; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130154.4]
  wire [5:0] _T_591; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130159.4]
  wire [12:0] real_hits; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130166.4]
  wire  _T_598; // @[TLB.scala 211:18:freechips.rocketchip.system.DefaultRV32Config.fir@130167.4]
  wire [13:0] hits; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130168.4]
  wire [33:0] _GEN_33; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130175.4]
  wire [33:0] _GEN_34; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130175.4]
  wire [33:0] _GEN_35; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130175.4]
  wire [33:0] _GEN_37; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130216.4]
  wire [33:0] _GEN_38; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130216.4]
  wire [33:0] _GEN_39; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130216.4]
  wire [33:0] _GEN_41; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130257.4]
  wire [33:0] _GEN_42; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130257.4]
  wire [33:0] _GEN_43; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130257.4]
  wire [33:0] _GEN_45; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130298.4]
  wire [33:0] _GEN_46; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130298.4]
  wire [33:0] _GEN_47; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130298.4]
  wire [33:0] _GEN_49; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130339.4]
  wire [33:0] _GEN_50; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130339.4]
  wire [33:0] _GEN_51; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130339.4]
  wire [33:0] _GEN_53; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130380.4]
  wire [33:0] _GEN_54; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130380.4]
  wire [33:0] _GEN_55; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130380.4]
  wire [33:0] _GEN_57; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130421.4]
  wire [33:0] _GEN_58; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130421.4]
  wire [33:0] _GEN_59; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130421.4]
  wire [33:0] _GEN_61; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130462.4]
  wire [33:0] _GEN_62; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130462.4]
  wire [33:0] _GEN_63; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130462.4]
  wire  _T_758; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@130527.4]
  wire [9:0] _T_761; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130538.4]
  wire [19:0] _T_765; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130542.4]
  wire [9:0] _T_766; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130543.4]
  wire [19:0] _T_767; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130544.4]
  wire  _T_782; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@130574.4]
  wire [9:0] _T_785; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130585.4]
  wire [19:0] _T_789; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130589.4]
  wire [9:0] _T_790; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130590.4]
  wire [19:0] _T_791; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130591.4]
  wire  _T_806; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@130621.4]
  wire [9:0] _T_809; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130632.4]
  wire [19:0] _T_813; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130636.4]
  wire [9:0] _T_814; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130637.4]
  wire [19:0] _T_815; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130638.4]
  wire  _T_830; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@130668.4]
  wire [9:0] _T_833; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130679.4]
  wire [19:0] _T_837; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130683.4]
  wire [9:0] _T_838; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130684.4]
  wire [19:0] _T_839; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130685.4]
  wire [9:0] _T_857; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130726.4]
  wire [19:0] _T_861; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130730.4]
  wire [9:0] _T_862; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130731.4]
  wire [19:0] _T_863; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130732.4]
  wire [19:0] _T_865; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130734.4]
  wire [19:0] _T_866; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130735.4]
  wire [19:0] _T_867; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130736.4]
  wire [19:0] _T_868; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130737.4]
  wire [19:0] _T_869; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130738.4]
  wire [19:0] _T_870; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130739.4]
  wire [19:0] _T_871; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130740.4]
  wire [19:0] _T_872; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130741.4]
  wire [19:0] _T_873; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130742.4]
  wire [19:0] _T_874; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130743.4]
  wire [19:0] _T_875; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130744.4]
  wire [19:0] _T_876; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130745.4]
  wire [19:0] _T_877; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130746.4]
  wire [19:0] _T_878; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130747.4]
  wire [19:0] _T_879; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130748.4]
  wire [19:0] _T_880; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130749.4]
  wire [19:0] _T_881; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130750.4]
  wire [19:0] _T_882; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130751.4]
  wire [19:0] _T_883; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130752.4]
  wire [19:0] _T_884; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130753.4]
  wire [19:0] _T_885; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130754.4]
  wire [19:0] _T_886; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130755.4]
  wire [19:0] _T_887; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130756.4]
  wire [19:0] _T_888; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130757.4]
  wire [19:0] _T_889; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130758.4]
  wire [19:0] _T_890; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130759.4]
  wire [19:0] ppn; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130760.4]
  wire  _T_892; // @[TLB.scala 215:22:freechips.rocketchip.system.DefaultRV32Config.fir@130763.4]
  wire  _T_893; // @[TLB.scala 215:19:freechips.rocketchip.system.DefaultRV32Config.fir@130764.4]
  wire  _T_895; // @[TLB.scala 221:25:freechips.rocketchip.system.DefaultRV32Config.fir@130771.6]
  wire  _T_896; // @[PTW.scala 68:47:freechips.rocketchip.system.DefaultRV32Config.fir@130774.6]
  wire  _T_897; // @[PTW.scala 68:44:freechips.rocketchip.system.DefaultRV32Config.fir@130775.6]
  wire  _T_898; // @[PTW.scala 68:38:freechips.rocketchip.system.DefaultRV32Config.fir@130776.6]
  wire  _T_899; // @[PTW.scala 68:32:freechips.rocketchip.system.DefaultRV32Config.fir@130777.6]
  wire  _T_900; // @[PTW.scala 68:52:freechips.rocketchip.system.DefaultRV32Config.fir@130778.6]
  wire  _T_901; // @[PTW.scala 72:35:freechips.rocketchip.system.DefaultRV32Config.fir@130779.6]
  wire  _T_907; // @[PTW.scala 73:35:freechips.rocketchip.system.DefaultRV32Config.fir@130786.6]
  wire  _T_908; // @[PTW.scala 73:40:freechips.rocketchip.system.DefaultRV32Config.fir@130787.6]
  wire  _T_914; // @[PTW.scala 74:35:freechips.rocketchip.system.DefaultRV32Config.fir@130794.6]
  wire  _T_915; // @[TLB.scala 234:37:freechips.rocketchip.system.DefaultRV32Config.fir@130803.6]
  wire [6:0] _T_923; // @[TLB.scala 136:26:freechips.rocketchip.system.DefaultRV32Config.fir@130815.8]
  wire [33:0] _T_931; // @[TLB.scala 136:26:freechips.rocketchip.system.DefaultRV32Config.fir@130823.8]
  wire  _T_932; // @[TLB.scala 236:40:freechips.rocketchip.system.DefaultRV32Config.fir@130827.8]
  wire  _T_933; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@130829.10]
  wire  _GEN_66; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@130830.10]
  wire  _T_948; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@130850.10]
  wire  _GEN_70; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@130851.10]
  wire  _T_963; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@130871.10]
  wire  _GEN_74; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@130872.10]
  wire  _T_978; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@130892.10]
  wire  _GEN_78; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@130893.10]
  wire [2:0] _T_993; // @[TLB.scala 241:22:freechips.rocketchip.system.DefaultRV32Config.fir@130915.10]
  wire  _T_994; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@130916.10]
  wire  _T_995; // @[TLB.scala 243:15:freechips.rocketchip.system.DefaultRV32Config.fir@130918.12]
  wire  _GEN_80; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130919.12]
  wire  _GEN_81; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130919.12]
  wire  _GEN_82; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130919.12]
  wire  _GEN_83; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130919.12]
  wire [1:0] _T_996; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@130927.12]
  wire  _GEN_950; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  wire  _GEN_84; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  wire  _GEN_951; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  wire  _GEN_85; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  wire  _GEN_952; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  wire  _GEN_86; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  wire  _GEN_953; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  wire  _GEN_87; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  wire  _GEN_92; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130917.10]
  wire  _GEN_93; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130917.10]
  wire  _GEN_94; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130917.10]
  wire  _GEN_95; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130917.10]
  wire  _T_1011; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@130945.10]
  wire  _GEN_102; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130948.12]
  wire  _GEN_103; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130948.12]
  wire  _GEN_104; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130948.12]
  wire  _GEN_105; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130948.12]
  wire  _GEN_106; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130957.12]
  wire  _GEN_107; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130957.12]
  wire  _GEN_108; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130957.12]
  wire  _GEN_109; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130957.12]
  wire  _GEN_114; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130946.10]
  wire  _GEN_115; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130946.10]
  wire  _GEN_116; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130946.10]
  wire  _GEN_117; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130946.10]
  wire  _T_1028; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@130974.10]
  wire  _GEN_124; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130977.12]
  wire  _GEN_125; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130977.12]
  wire  _GEN_126; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130977.12]
  wire  _GEN_127; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130977.12]
  wire  _GEN_128; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130986.12]
  wire  _GEN_129; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130986.12]
  wire  _GEN_130; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130986.12]
  wire  _GEN_131; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130986.12]
  wire  _GEN_136; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130975.10]
  wire  _GEN_137; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130975.10]
  wire  _GEN_138; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130975.10]
  wire  _GEN_139; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130975.10]
  wire  _T_1045; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131003.10]
  wire  _GEN_146; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131006.12]
  wire  _GEN_147; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131006.12]
  wire  _GEN_148; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131006.12]
  wire  _GEN_149; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131006.12]
  wire  _GEN_150; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131015.12]
  wire  _GEN_151; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131015.12]
  wire  _GEN_152; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131015.12]
  wire  _GEN_153; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131015.12]
  wire  _GEN_158; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131004.10]
  wire  _GEN_159; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131004.10]
  wire  _GEN_160; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131004.10]
  wire  _GEN_161; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131004.10]
  wire  _T_1062; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131032.10]
  wire  _GEN_168; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131035.12]
  wire  _GEN_169; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131035.12]
  wire  _GEN_170; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131035.12]
  wire  _GEN_171; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131035.12]
  wire  _GEN_172; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131044.12]
  wire  _GEN_173; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131044.12]
  wire  _GEN_174; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131044.12]
  wire  _GEN_175; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131044.12]
  wire  _GEN_180; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131033.10]
  wire  _GEN_181; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131033.10]
  wire  _GEN_182; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131033.10]
  wire  _GEN_183; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131033.10]
  wire  _T_1079; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131061.10]
  wire  _GEN_190; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131064.12]
  wire  _GEN_191; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131064.12]
  wire  _GEN_192; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131064.12]
  wire  _GEN_193; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131064.12]
  wire  _GEN_194; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131073.12]
  wire  _GEN_195; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131073.12]
  wire  _GEN_196; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131073.12]
  wire  _GEN_197; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131073.12]
  wire  _GEN_202; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131062.10]
  wire  _GEN_203; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131062.10]
  wire  _GEN_204; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131062.10]
  wire  _GEN_205; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131062.10]
  wire  _T_1096; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131090.10]
  wire  _GEN_212; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131093.12]
  wire  _GEN_213; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131093.12]
  wire  _GEN_214; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131093.12]
  wire  _GEN_215; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131093.12]
  wire  _GEN_216; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131102.12]
  wire  _GEN_217; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131102.12]
  wire  _GEN_218; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131102.12]
  wire  _GEN_219; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131102.12]
  wire  _GEN_224; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131091.10]
  wire  _GEN_225; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131091.10]
  wire  _GEN_226; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131091.10]
  wire  _GEN_227; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131091.10]
  wire  _T_1113; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131119.10]
  wire  _GEN_234; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131122.12]
  wire  _GEN_235; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131122.12]
  wire  _GEN_236; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131122.12]
  wire  _GEN_237; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131122.12]
  wire  _GEN_238; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131131.12]
  wire  _GEN_239; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131131.12]
  wire  _GEN_240; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131131.12]
  wire  _GEN_241; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131131.12]
  wire  _GEN_246; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131120.10]
  wire  _GEN_247; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131120.10]
  wire  _GEN_248; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131120.10]
  wire  _GEN_249; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131120.10]
  wire  _GEN_258; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_262; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_266; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_270; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_272; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_273; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_274; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_275; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_282; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_283; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_284; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_285; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_292; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_293; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_294; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_295; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_302; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_303; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_304; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_305; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_312; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_313; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_314; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_315; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_322; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_323; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_324; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_325; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_332; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_333; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_334; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_335; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_342; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_343; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_344; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_345; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  wire  _GEN_354; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_358; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_362; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_366; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_370; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_372; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_373; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_374; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_375; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_382; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_383; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_384; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_385; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_392; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_393; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_394; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_395; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_402; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_403; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_404; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_405; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_412; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_413; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_414; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_415; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_422; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_423; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_424; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_425; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_432; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_433; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_434; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_435; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_442; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_443; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_444; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_445; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  wire  _GEN_454; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_458; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_462; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_466; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_470; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_472; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_473; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_474; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_475; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_482; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_483; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_484; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_485; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_492; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_493; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_494; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_495; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_502; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_503; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_504; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_505; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_512; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_513; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_514; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_515; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_522; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_523; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_524; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_525; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_532; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_533; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_534; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_535; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_542; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_543; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_544; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire  _GEN_545; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  wire [5:0] _T_1575; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132170.4]
  wire [13:0] ptw_ae_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132178.4]
  wire [5:0] _T_1589; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132185.4]
  wire [12:0] _T_1596; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132192.4]
  wire [12:0] _T_1610; // @[TLB.scala 253:98:freechips.rocketchip.system.DefaultRV32Config.fir@132206.4]
  wire [12:0] priv_x_ok; // @[TLB.scala 254:22:freechips.rocketchip.system.DefaultRV32Config.fir@132234.4]
  wire [5:0] _T_1653; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132251.4]
  wire [12:0] _T_1660; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132258.4]
  wire [12:0] _T_1689; // @[TLB.scala 257:39:freechips.rocketchip.system.DefaultRV32Config.fir@132289.4]
  wire [13:0] x_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132290.4]
  wire [13:0] _T_1704; // @[TLB.scala 258:89:freechips.rocketchip.system.DefaultRV32Config.fir@132305.4]
  wire [1:0] _T_1721; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@132324.4]
  wire [5:0] _T_1726; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132329.4]
  wire [13:0] _T_1733; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132336.4]
  wire [13:0] px_array; // @[TLB.scala 260:87:freechips.rocketchip.system.DefaultRV32Config.fir@132338.4]
  wire [1:0] _T_1749; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@132354.4]
  wire [5:0] _T_1754; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132359.4]
  wire [13:0] c_array; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132366.4]
  wire [13:0] _T_1900; // @[TLB.scala 305:33:freechips.rocketchip.system.DefaultRV32Config.fir@132527.4]
  wire [13:0] pf_inst_array; // @[TLB.scala 305:23:freechips.rocketchip.system.DefaultRV32Config.fir@132528.4]
  wire  tlb_hit; // @[TLB.scala 307:27:freechips.rocketchip.system.DefaultRV32Config.fir@132529.4]
  wire  _T_1903; // @[TLB.scala 308:43:freechips.rocketchip.system.DefaultRV32Config.fir@132532.4]
  wire  tlb_miss; // @[TLB.scala 308:40:freechips.rocketchip.system.DefaultRV32Config.fir@132533.4]
  reg [6:0] _T_1904; // @[Replacement.scala 41:30:freechips.rocketchip.system.DefaultRV32Config.fir@132534.4]
  reg [31:0] _RAND_94;
  reg [2:0] _T_1905; // @[Replacement.scala 41:30:freechips.rocketchip.system.DefaultRV32Config.fir@132535.4]
  reg [31:0] _RAND_95;
  wire  _T_1906; // @[TLB.scala 312:22:freechips.rocketchip.system.DefaultRV32Config.fir@132536.4]
  wire  _T_1907; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132538.6]
  wire  _T_1908; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132539.6]
  wire  _T_1909; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132540.6]
  wire  _T_1910; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132541.6]
  wire  _T_1911; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132542.6]
  wire  _T_1912; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132543.6]
  wire  _T_1913; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132544.6]
  wire [7:0] _T_1920; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132552.8]
  wire [3:0] _T_1921; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@132553.8]
  wire [3:0] _T_1922; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@132554.8]
  wire  _T_1923; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@132555.8]
  wire [3:0] _T_1924; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@132556.8]
  wire [1:0] _T_1925; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@132557.8]
  wire [1:0] _T_1926; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@132558.8]
  wire  _T_1927; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@132559.8]
  wire [1:0] _T_1928; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@132560.8]
  wire  _T_1929; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@132561.8]
  wire [2:0] _T_1931; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132563.8]
  wire [7:0] _T_1932; // @[Replacement.scala 46:28:freechips.rocketchip.system.DefaultRV32Config.fir@132564.8]
  wire  _T_1933; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132565.8]
  wire  _T_1934; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132566.8]
  wire [7:0] _T_1936; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132568.8]
  wire [7:0] _T_1937; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132569.8]
  wire [7:0] _T_1938; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132570.8]
  wire [7:0] _T_1939; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132571.8]
  wire [7:0] _T_1940; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132572.8]
  wire [1:0] _T_1941; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132573.8]
  wire  _T_1942; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132574.8]
  wire  _T_1943; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132575.8]
  wire [3:0] _T_1944; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132576.8]
  wire [7:0] _GEN_983; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132577.8]
  wire [7:0] _T_1945; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132577.8]
  wire [7:0] _T_1946; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132578.8]
  wire [7:0] _T_1947; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132579.8]
  wire [7:0] _T_1948; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132580.8]
  wire [7:0] _T_1949; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132581.8]
  wire [2:0] _T_1950; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132582.8]
  wire  _T_1951; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132583.8]
  wire  _T_1952; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132584.8]
  wire [7:0] _T_1953; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132585.8]
  wire [7:0] _T_1954; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132586.8]
  wire [7:0] _T_1955; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132587.8]
  wire [7:0] _T_1956; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132588.8]
  wire [7:0] _T_1957; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132589.8]
  wire [7:0] _T_1958; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132590.8]
  wire [6:0] _T_1960; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@132592.8]
  wire  _T_1961; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132595.6]
  wire  _T_1962; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132596.6]
  wire  _T_1963; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132597.6]
  wire [3:0] _T_1966; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132601.8]
  wire [1:0] _T_1967; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@132602.8]
  wire [1:0] _T_1968; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@132603.8]
  wire  _T_1969; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@132604.8]
  wire [1:0] _T_1970; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@132605.8]
  wire  _T_1971; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@132606.8]
  wire [1:0] _T_1972; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132607.8]
  wire [3:0] _T_1973; // @[Replacement.scala 46:28:freechips.rocketchip.system.DefaultRV32Config.fir@132608.8]
  wire  _T_1974; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132609.8]
  wire  _T_1975; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132610.8]
  wire [3:0] _T_1977; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132612.8]
  wire [3:0] _T_1978; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132613.8]
  wire [3:0] _T_1979; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132614.8]
  wire [3:0] _T_1980; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132615.8]
  wire [3:0] _T_1981; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132616.8]
  wire [1:0] _T_1982; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132617.8]
  wire  _T_1983; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132618.8]
  wire  _T_1984; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132619.8]
  wire [3:0] _T_1985; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132620.8]
  wire [3:0] _T_1986; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132621.8]
  wire [3:0] _T_1987; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132622.8]
  wire [3:0] _T_1988; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132623.8]
  wire [3:0] _T_1989; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132624.8]
  wire [3:0] _T_1990; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132625.8]
  wire [2:0] _T_1992; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@132627.8]
  wire [5:0] _T_1993; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132631.4]
  wire [2:0] _T_1994; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132632.4]
  wire  _T_1995; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132633.4]
  wire [1:0] _T_1997; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132635.4]
  wire  _T_1998; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132636.4]
  wire  _T_2000; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132638.4]
  wire  _T_2002; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132640.4]
  wire  _T_2004; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132642.4]
  wire  _T_2006; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132644.4]
  wire  _T_2008; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132646.4]
  wire  _T_2009; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132647.4]
  wire [2:0] _T_2010; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132648.4]
  wire  _T_2011; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132649.4]
  wire [1:0] _T_2013; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132651.4]
  wire  _T_2014; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132652.4]
  wire  _T_2016; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132654.4]
  wire  _T_2018; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132656.4]
  wire  _T_2020; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132658.4]
  wire  _T_2022; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132660.4]
  wire  _T_2024; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132662.4]
  wire  _T_2025; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132663.4]
  wire  _T_2026; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132664.4]
  wire  _T_2027; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@132665.4]
  wire  _T_2028; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132666.4]
  wire  _T_2029; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132667.4]
  wire [6:0] _T_2030; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132668.4]
  wire [2:0] _T_2031; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132669.4]
  wire  _T_2032; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132670.4]
  wire [1:0] _T_2034; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132672.4]
  wire  _T_2035; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132673.4]
  wire  _T_2037; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132675.4]
  wire  _T_2039; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132677.4]
  wire  _T_2041; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132679.4]
  wire  _T_2043; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132681.4]
  wire  _T_2045; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132683.4]
  wire  _T_2046; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132684.4]
  wire [3:0] _T_2047; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132685.4]
  wire [1:0] _T_2048; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132686.4]
  wire  _T_2049; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132687.4]
  wire  _T_2051; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132689.4]
  wire  _T_2053; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132691.4]
  wire  _T_2055; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132693.4]
  wire [1:0] _T_2057; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132695.4]
  wire  _T_2058; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132696.4]
  wire  _T_2060; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132698.4]
  wire  _T_2062; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132700.4]
  wire  _T_2064; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132702.4]
  wire  _T_2066; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132704.4]
  wire  _T_2067; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@132705.4]
  wire  _T_2068; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132706.4]
  wire  _T_2069; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132707.4]
  wire  _T_2070; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132708.4]
  wire  _T_2071; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@132709.4]
  wire  _T_2072; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132710.4]
  wire  _T_2073; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132711.4]
  wire  _T_2075; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@132713.4]
  wire  _T_2076; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132714.4]
  wire  multipleHits; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132715.4]
  wire [13:0] _T_2086; // @[TLB.scala 327:47:freechips.rocketchip.system.DefaultRV32Config.fir@132728.4]
  wire [13:0] _T_2093; // @[TLB.scala 330:23:freechips.rocketchip.system.DefaultRV32Config.fir@132738.4]
  wire [13:0] _T_2094; // @[TLB.scala 330:33:freechips.rocketchip.system.DefaultRV32Config.fir@132739.4]
  wire [13:0] _T_2100; // @[TLB.scala 334:33:freechips.rocketchip.system.DefaultRV32Config.fir@132749.4]
  wire  _T_2107; // @[TLB.scala 337:29:freechips.rocketchip.system.DefaultRV32Config.fir@132759.4]
  wire  _T_2113; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@132770.4]
  wire  _T_2114; // @[TLB.scala 346:25:freechips.rocketchip.system.DefaultRV32Config.fir@132771.4]
  wire [2:0] _GEN_985; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132779.6]
  wire [3:0] _T_2119; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132779.6]
  wire  _T_2120; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132780.6]
  wire [1:0] _T_2122; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132782.6]
  wire [3:0] _T_2126; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132786.6]
  wire  _T_2127; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132787.6]
  wire [2:0] _T_2129; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132789.6]
  wire [1:0] _T_2130; // @[Replacement.scala 63:8:freechips.rocketchip.system.DefaultRV32Config.fir@132790.6]
  wire [3:0] _T_2133; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132793.6]
  wire  _T_2134; // @[TLB.scala 394:16:freechips.rocketchip.system.DefaultRV32Config.fir@132794.6]
  wire [3:0] _T_2135; // @[TLB.scala 394:43:freechips.rocketchip.system.DefaultRV32Config.fir@132795.6]
  wire  _T_2136; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132796.6]
  wire  _T_2137; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132797.6]
  wire  _T_2138; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132798.6]
  wire [6:0] _GEN_986; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132809.6]
  wire [7:0] _T_2148; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132809.6]
  wire  _T_2149; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132810.6]
  wire [1:0] _T_2151; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132812.6]
  wire [7:0] _T_2155; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132816.6]
  wire  _T_2156; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132817.6]
  wire [2:0] _T_2158; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132819.6]
  wire [7:0] _T_2162; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132823.6]
  wire  _T_2163; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132824.6]
  wire [3:0] _T_2165; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132826.6]
  wire [2:0] _T_2166; // @[Replacement.scala 63:8:freechips.rocketchip.system.DefaultRV32Config.fir@132827.6]
  wire [7:0] _T_2197; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132858.6]
  wire  _T_2198; // @[TLB.scala 394:16:freechips.rocketchip.system.DefaultRV32Config.fir@132859.6]
  wire [7:0] _T_2199; // @[TLB.scala 394:43:freechips.rocketchip.system.DefaultRV32Config.fir@132860.6]
  wire  _T_2200; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132861.6]
  wire  _T_2201; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132862.6]
  wire  _T_2202; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132863.6]
  wire  _T_2203; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132864.6]
  wire  _T_2204; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132865.6]
  wire  _T_2205; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132866.6]
  wire  _T_2206; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132867.6]
  wire  _T_2243; // @[TLB.scala 360:17:freechips.rocketchip.system.DefaultRV32Config.fir@132919.4]
  wire  _T_2244; // @[TLB.scala 360:28:freechips.rocketchip.system.DefaultRV32Config.fir@132920.4]
  wire  _T_2245; // @[TLB.scala 368:14:freechips.rocketchip.system.DefaultRV32Config.fir@132928.6]
  wire [19:0] _T_2246; // @[TLB.scala 368:58:freechips.rocketchip.system.DefaultRV32Config.fir@132929.6]
  wire  _T_2247; // @[TLB.scala 368:72:freechips.rocketchip.system.DefaultRV32Config.fir@132930.6]
  wire  _T_2248; // @[TLB.scala 368:34:freechips.rocketchip.system.DefaultRV32Config.fir@132931.6]
  wire  _T_2250; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@132933.6]
  wire  _T_2251; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@132934.6]
  wire [9:0] _T_2257; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@132948.8]
  wire  _T_2258; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@132949.8]
  wire  _T_2261; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@132956.10]
  wire  _T_2273; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@132980.10]
  wire  _T_2278; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@132991.10]
  wire  _T_2290; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133015.10]
  wire  _T_2295; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133026.10]
  wire  _T_2307; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133050.10]
  wire  _T_2312; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133061.10]
  wire  _T_2324; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133085.10]
  wire  _T_2395; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133247.10]
  wire  _GEN_648; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133248.10]
  wire  _T_2396; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133251.10]
  wire  _GEN_649; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133252.10]
  wire  _T_2397; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133255.10]
  wire  _GEN_650; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133256.10]
  wire  _T_2398; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133259.10]
  wire  _GEN_651; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133260.10]
  wire  _GEN_652; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133106.8]
  wire  _GEN_653; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133106.8]
  wire  _GEN_654; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133106.8]
  wire  _GEN_655; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133106.8]
  wire [9:0] _T_2404; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@133279.8]
  wire  _T_2405; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@133280.8]
  wire  _T_2408; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133287.10]
  wire  _T_2420; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133311.10]
  wire  _T_2425; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133322.10]
  wire  _T_2437; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133346.10]
  wire  _T_2442; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133357.10]
  wire  _T_2454; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133381.10]
  wire  _T_2459; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133392.10]
  wire  _T_2471; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133416.10]
  wire  _T_2542; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133578.10]
  wire  _GEN_676; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133579.10]
  wire  _T_2543; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133582.10]
  wire  _GEN_677; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133583.10]
  wire  _T_2544; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133586.10]
  wire  _GEN_678; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133587.10]
  wire  _T_2545; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133590.10]
  wire  _GEN_679; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133591.10]
  wire  _GEN_680; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133437.8]
  wire  _GEN_681; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133437.8]
  wire  _GEN_682; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133437.8]
  wire  _GEN_683; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133437.8]
  wire [9:0] _T_2551; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@133610.8]
  wire  _T_2552; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@133611.8]
  wire  _T_2555; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133618.10]
  wire  _T_2567; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133642.10]
  wire  _T_2572; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133653.10]
  wire  _T_2584; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133677.10]
  wire  _T_2589; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133688.10]
  wire  _T_2601; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133712.10]
  wire  _T_2606; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133723.10]
  wire  _T_2618; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133747.10]
  wire  _T_2689; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133909.10]
  wire  _GEN_704; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133910.10]
  wire  _T_2690; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133913.10]
  wire  _GEN_705; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133914.10]
  wire  _T_2691; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133917.10]
  wire  _GEN_706; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133918.10]
  wire  _T_2692; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133921.10]
  wire  _GEN_707; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133922.10]
  wire  _GEN_708; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133768.8]
  wire  _GEN_709; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133768.8]
  wire  _GEN_710; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133768.8]
  wire  _GEN_711; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133768.8]
  wire [9:0] _T_2698; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@133941.8]
  wire  _T_2699; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@133942.8]
  wire  _T_2702; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133949.10]
  wire  _T_2714; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133973.10]
  wire  _T_2719; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133984.10]
  wire  _T_2731; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134008.10]
  wire  _T_2736; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134019.10]
  wire  _T_2748; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134043.10]
  wire  _T_2753; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134054.10]
  wire  _T_2765; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134078.10]
  wire  _T_2836; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134240.10]
  wire  _GEN_732; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134241.10]
  wire  _T_2837; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134244.10]
  wire  _GEN_733; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134245.10]
  wire  _T_2838; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134248.10]
  wire  _GEN_734; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134249.10]
  wire  _T_2839; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134252.10]
  wire  _GEN_735; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134253.10]
  wire  _GEN_736; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134099.8]
  wire  _GEN_737; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134099.8]
  wire  _GEN_738; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134099.8]
  wire  _GEN_739; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134099.8]
  wire [9:0] _T_2845; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@134272.8]
  wire  _T_2846; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@134273.8]
  wire  _T_2849; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134280.10]
  wire  _T_2861; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134304.10]
  wire  _T_2866; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134315.10]
  wire  _T_2878; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134339.10]
  wire  _T_2883; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134350.10]
  wire  _T_2895; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134374.10]
  wire  _T_2900; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134385.10]
  wire  _T_2912; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134409.10]
  wire  _T_2983; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134571.10]
  wire  _GEN_760; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134572.10]
  wire  _T_2984; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134575.10]
  wire  _GEN_761; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134576.10]
  wire  _T_2985; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134579.10]
  wire  _GEN_762; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134580.10]
  wire  _T_2986; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134583.10]
  wire  _GEN_763; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134584.10]
  wire  _GEN_764; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134430.8]
  wire  _GEN_765; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134430.8]
  wire  _GEN_766; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134430.8]
  wire  _GEN_767; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134430.8]
  wire [9:0] _T_2992; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@134603.8]
  wire  _T_2993; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@134604.8]
  wire  _T_2996; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134611.10]
  wire  _T_3008; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134635.10]
  wire  _T_3013; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134646.10]
  wire  _T_3025; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134670.10]
  wire  _T_3030; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134681.10]
  wire  _T_3042; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134705.10]
  wire  _T_3047; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134716.10]
  wire  _T_3059; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134740.10]
  wire  _T_3130; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134902.10]
  wire  _GEN_788; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134903.10]
  wire  _T_3131; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134906.10]
  wire  _GEN_789; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134907.10]
  wire  _T_3132; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134910.10]
  wire  _GEN_790; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134911.10]
  wire  _T_3133; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134914.10]
  wire  _GEN_791; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134915.10]
  wire  _GEN_792; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134761.8]
  wire  _GEN_793; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134761.8]
  wire  _GEN_794; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134761.8]
  wire  _GEN_795; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134761.8]
  wire [9:0] _T_3139; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@134934.8]
  wire  _T_3140; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@134935.8]
  wire  _T_3143; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134942.10]
  wire  _T_3155; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134966.10]
  wire  _T_3160; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134977.10]
  wire  _T_3172; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135001.10]
  wire  _T_3177; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135012.10]
  wire  _T_3189; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135036.10]
  wire  _T_3194; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135047.10]
  wire  _T_3206; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135071.10]
  wire  _T_3277; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135233.10]
  wire  _GEN_816; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135234.10]
  wire  _T_3278; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135237.10]
  wire  _GEN_817; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135238.10]
  wire  _T_3279; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135241.10]
  wire  _GEN_818; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135242.10]
  wire  _T_3280; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135245.10]
  wire  _GEN_819; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135246.10]
  wire  _GEN_820; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135092.8]
  wire  _GEN_821; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135092.8]
  wire  _GEN_822; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135092.8]
  wire  _GEN_823; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135092.8]
  wire [9:0] _T_3286; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@135265.8]
  wire  _T_3287; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@135266.8]
  wire  _T_3290; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135273.10]
  wire  _T_3302; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135297.10]
  wire  _T_3307; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135308.10]
  wire  _T_3319; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135332.10]
  wire  _T_3324; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135343.10]
  wire  _T_3336; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135367.10]
  wire  _T_3341; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135378.10]
  wire  _T_3353; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135402.10]
  wire  _T_3424; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135564.10]
  wire  _GEN_844; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135565.10]
  wire  _T_3425; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135568.10]
  wire  _GEN_845; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135569.10]
  wire  _T_3426; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135572.10]
  wire  _GEN_846; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135573.10]
  wire  _T_3427; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135576.10]
  wire  _GEN_847; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135577.10]
  wire  _GEN_848; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135423.8]
  wire  _GEN_849; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135423.8]
  wire  _GEN_850; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135423.8]
  wire  _GEN_851; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135423.8]
  wire  _T_3459; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135643.10]
  wire  _GEN_857; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135644.10]
  wire  _GEN_858; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135607.8]
  wire  _T_3491; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135707.10]
  wire  _GEN_861; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135708.10]
  wire  _GEN_862; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135671.8]
  wire  _T_3523; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135771.10]
  wire  _GEN_865; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135772.10]
  wire  _GEN_866; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135735.8]
  wire  _T_3555; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135835.10]
  wire  _GEN_869; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135836.10]
  wire  _GEN_870; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135799.8]
  wire  _T_3587; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135899.10]
  wire  _GEN_873; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135900.10]
  wire  _GEN_874; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135863.8]
  wire  _T_3589; // @[TLB.scala 375:24:freechips.rocketchip.system.DefaultRV32Config.fir@135909.4]
  _2_1 _2 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@129520.4]
    .io_x_ppn(_2_io_x_ppn),
    .io_x_u(_2_io_x_u),
    .io_x_ae(_2_io_x_ae),
    .io_x_sw(_2_io_x_sw),
    .io_x_sx(_2_io_x_sx),
    .io_x_sr(_2_io_x_sr),
    .io_x_pw(_2_io_x_pw),
    .io_x_px(_2_io_x_px),
    .io_x_pr(_2_io_x_pr),
    .io_x_pal(_2_io_x_pal),
    .io_x_paa(_2_io_x_paa),
    .io_x_eff(_2_io_x_eff),
    .io_x_c(_2_io_x_c),
    .io_y_ppn(_2_io_y_ppn),
    .io_y_u(_2_io_y_u),
    .io_y_ae(_2_io_y_ae),
    .io_y_sw(_2_io_y_sw),
    .io_y_sx(_2_io_y_sx),
    .io_y_sr(_2_io_y_sr),
    .io_y_pw(_2_io_y_pw),
    .io_y_px(_2_io_y_px),
    .io_y_pr(_2_io_y_pr),
    .io_y_pal(_2_io_y_pal),
    .io_y_paa(_2_io_y_paa),
    .io_y_eff(_2_io_y_eff),
    .io_y_c(_2_io_y_c)
  );
  PMPChecker pmp ( // @[TLB.scala 189:19:freechips.rocketchip.system.DefaultRV32Config.fir@129541.4]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x)
  );
  _2_1 _2_1 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130206.4]
    .io_x_ppn(_2_1_io_x_ppn),
    .io_x_u(_2_1_io_x_u),
    .io_x_ae(_2_1_io_x_ae),
    .io_x_sw(_2_1_io_x_sw),
    .io_x_sx(_2_1_io_x_sx),
    .io_x_sr(_2_1_io_x_sr),
    .io_x_pw(_2_1_io_x_pw),
    .io_x_px(_2_1_io_x_px),
    .io_x_pr(_2_1_io_x_pr),
    .io_x_pal(_2_1_io_x_pal),
    .io_x_paa(_2_1_io_x_paa),
    .io_x_eff(_2_1_io_x_eff),
    .io_x_c(_2_1_io_x_c),
    .io_y_ppn(_2_1_io_y_ppn),
    .io_y_u(_2_1_io_y_u),
    .io_y_ae(_2_1_io_y_ae),
    .io_y_sw(_2_1_io_y_sw),
    .io_y_sx(_2_1_io_y_sx),
    .io_y_sr(_2_1_io_y_sr),
    .io_y_pw(_2_1_io_y_pw),
    .io_y_px(_2_1_io_y_px),
    .io_y_pr(_2_1_io_y_pr),
    .io_y_pal(_2_1_io_y_pal),
    .io_y_paa(_2_1_io_y_paa),
    .io_y_eff(_2_1_io_y_eff),
    .io_y_c(_2_1_io_y_c)
  );
  _2_1 _2_2 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130247.4]
    .io_x_ppn(_2_2_io_x_ppn),
    .io_x_u(_2_2_io_x_u),
    .io_x_ae(_2_2_io_x_ae),
    .io_x_sw(_2_2_io_x_sw),
    .io_x_sx(_2_2_io_x_sx),
    .io_x_sr(_2_2_io_x_sr),
    .io_x_pw(_2_2_io_x_pw),
    .io_x_px(_2_2_io_x_px),
    .io_x_pr(_2_2_io_x_pr),
    .io_x_pal(_2_2_io_x_pal),
    .io_x_paa(_2_2_io_x_paa),
    .io_x_eff(_2_2_io_x_eff),
    .io_x_c(_2_2_io_x_c),
    .io_y_ppn(_2_2_io_y_ppn),
    .io_y_u(_2_2_io_y_u),
    .io_y_ae(_2_2_io_y_ae),
    .io_y_sw(_2_2_io_y_sw),
    .io_y_sx(_2_2_io_y_sx),
    .io_y_sr(_2_2_io_y_sr),
    .io_y_pw(_2_2_io_y_pw),
    .io_y_px(_2_2_io_y_px),
    .io_y_pr(_2_2_io_y_pr),
    .io_y_pal(_2_2_io_y_pal),
    .io_y_paa(_2_2_io_y_paa),
    .io_y_eff(_2_2_io_y_eff),
    .io_y_c(_2_2_io_y_c)
  );
  _2_1 _2_3 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130288.4]
    .io_x_ppn(_2_3_io_x_ppn),
    .io_x_u(_2_3_io_x_u),
    .io_x_ae(_2_3_io_x_ae),
    .io_x_sw(_2_3_io_x_sw),
    .io_x_sx(_2_3_io_x_sx),
    .io_x_sr(_2_3_io_x_sr),
    .io_x_pw(_2_3_io_x_pw),
    .io_x_px(_2_3_io_x_px),
    .io_x_pr(_2_3_io_x_pr),
    .io_x_pal(_2_3_io_x_pal),
    .io_x_paa(_2_3_io_x_paa),
    .io_x_eff(_2_3_io_x_eff),
    .io_x_c(_2_3_io_x_c),
    .io_y_ppn(_2_3_io_y_ppn),
    .io_y_u(_2_3_io_y_u),
    .io_y_ae(_2_3_io_y_ae),
    .io_y_sw(_2_3_io_y_sw),
    .io_y_sx(_2_3_io_y_sx),
    .io_y_sr(_2_3_io_y_sr),
    .io_y_pw(_2_3_io_y_pw),
    .io_y_px(_2_3_io_y_px),
    .io_y_pr(_2_3_io_y_pr),
    .io_y_pal(_2_3_io_y_pal),
    .io_y_paa(_2_3_io_y_paa),
    .io_y_eff(_2_3_io_y_eff),
    .io_y_c(_2_3_io_y_c)
  );
  _2_1 _2_4 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130329.4]
    .io_x_ppn(_2_4_io_x_ppn),
    .io_x_u(_2_4_io_x_u),
    .io_x_ae(_2_4_io_x_ae),
    .io_x_sw(_2_4_io_x_sw),
    .io_x_sx(_2_4_io_x_sx),
    .io_x_sr(_2_4_io_x_sr),
    .io_x_pw(_2_4_io_x_pw),
    .io_x_px(_2_4_io_x_px),
    .io_x_pr(_2_4_io_x_pr),
    .io_x_pal(_2_4_io_x_pal),
    .io_x_paa(_2_4_io_x_paa),
    .io_x_eff(_2_4_io_x_eff),
    .io_x_c(_2_4_io_x_c),
    .io_y_ppn(_2_4_io_y_ppn),
    .io_y_u(_2_4_io_y_u),
    .io_y_ae(_2_4_io_y_ae),
    .io_y_sw(_2_4_io_y_sw),
    .io_y_sx(_2_4_io_y_sx),
    .io_y_sr(_2_4_io_y_sr),
    .io_y_pw(_2_4_io_y_pw),
    .io_y_px(_2_4_io_y_px),
    .io_y_pr(_2_4_io_y_pr),
    .io_y_pal(_2_4_io_y_pal),
    .io_y_paa(_2_4_io_y_paa),
    .io_y_eff(_2_4_io_y_eff),
    .io_y_c(_2_4_io_y_c)
  );
  _2_1 _2_5 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130370.4]
    .io_x_ppn(_2_5_io_x_ppn),
    .io_x_u(_2_5_io_x_u),
    .io_x_ae(_2_5_io_x_ae),
    .io_x_sw(_2_5_io_x_sw),
    .io_x_sx(_2_5_io_x_sx),
    .io_x_sr(_2_5_io_x_sr),
    .io_x_pw(_2_5_io_x_pw),
    .io_x_px(_2_5_io_x_px),
    .io_x_pr(_2_5_io_x_pr),
    .io_x_pal(_2_5_io_x_pal),
    .io_x_paa(_2_5_io_x_paa),
    .io_x_eff(_2_5_io_x_eff),
    .io_x_c(_2_5_io_x_c),
    .io_y_ppn(_2_5_io_y_ppn),
    .io_y_u(_2_5_io_y_u),
    .io_y_ae(_2_5_io_y_ae),
    .io_y_sw(_2_5_io_y_sw),
    .io_y_sx(_2_5_io_y_sx),
    .io_y_sr(_2_5_io_y_sr),
    .io_y_pw(_2_5_io_y_pw),
    .io_y_px(_2_5_io_y_px),
    .io_y_pr(_2_5_io_y_pr),
    .io_y_pal(_2_5_io_y_pal),
    .io_y_paa(_2_5_io_y_paa),
    .io_y_eff(_2_5_io_y_eff),
    .io_y_c(_2_5_io_y_c)
  );
  _2_1 _2_6 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130411.4]
    .io_x_ppn(_2_6_io_x_ppn),
    .io_x_u(_2_6_io_x_u),
    .io_x_ae(_2_6_io_x_ae),
    .io_x_sw(_2_6_io_x_sw),
    .io_x_sx(_2_6_io_x_sx),
    .io_x_sr(_2_6_io_x_sr),
    .io_x_pw(_2_6_io_x_pw),
    .io_x_px(_2_6_io_x_px),
    .io_x_pr(_2_6_io_x_pr),
    .io_x_pal(_2_6_io_x_pal),
    .io_x_paa(_2_6_io_x_paa),
    .io_x_eff(_2_6_io_x_eff),
    .io_x_c(_2_6_io_x_c),
    .io_y_ppn(_2_6_io_y_ppn),
    .io_y_u(_2_6_io_y_u),
    .io_y_ae(_2_6_io_y_ae),
    .io_y_sw(_2_6_io_y_sw),
    .io_y_sx(_2_6_io_y_sx),
    .io_y_sr(_2_6_io_y_sr),
    .io_y_pw(_2_6_io_y_pw),
    .io_y_px(_2_6_io_y_px),
    .io_y_pr(_2_6_io_y_pr),
    .io_y_pal(_2_6_io_y_pal),
    .io_y_paa(_2_6_io_y_paa),
    .io_y_eff(_2_6_io_y_eff),
    .io_y_c(_2_6_io_y_c)
  );
  _2_1 _2_7 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130452.4]
    .io_x_ppn(_2_7_io_x_ppn),
    .io_x_u(_2_7_io_x_u),
    .io_x_ae(_2_7_io_x_ae),
    .io_x_sw(_2_7_io_x_sw),
    .io_x_sx(_2_7_io_x_sx),
    .io_x_sr(_2_7_io_x_sr),
    .io_x_pw(_2_7_io_x_pw),
    .io_x_px(_2_7_io_x_px),
    .io_x_pr(_2_7_io_x_pr),
    .io_x_pal(_2_7_io_x_pal),
    .io_x_paa(_2_7_io_x_paa),
    .io_x_eff(_2_7_io_x_eff),
    .io_x_c(_2_7_io_x_c),
    .io_y_ppn(_2_7_io_y_ppn),
    .io_y_u(_2_7_io_y_u),
    .io_y_ae(_2_7_io_y_ae),
    .io_y_sw(_2_7_io_y_sw),
    .io_y_sx(_2_7_io_y_sx),
    .io_y_sr(_2_7_io_y_sr),
    .io_y_pw(_2_7_io_y_pw),
    .io_y_px(_2_7_io_y_px),
    .io_y_pr(_2_7_io_y_pr),
    .io_y_pal(_2_7_io_y_pal),
    .io_y_paa(_2_7_io_y_paa),
    .io_y_eff(_2_7_io_y_eff),
    .io_y_c(_2_7_io_y_c)
  );
  _2_1 _2_8 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130493.4]
    .io_x_ppn(_2_8_io_x_ppn),
    .io_x_u(_2_8_io_x_u),
    .io_x_ae(_2_8_io_x_ae),
    .io_x_sw(_2_8_io_x_sw),
    .io_x_sx(_2_8_io_x_sx),
    .io_x_sr(_2_8_io_x_sr),
    .io_x_pw(_2_8_io_x_pw),
    .io_x_px(_2_8_io_x_px),
    .io_x_pr(_2_8_io_x_pr),
    .io_x_pal(_2_8_io_x_pal),
    .io_x_paa(_2_8_io_x_paa),
    .io_x_eff(_2_8_io_x_eff),
    .io_x_c(_2_8_io_x_c),
    .io_y_ppn(_2_8_io_y_ppn),
    .io_y_u(_2_8_io_y_u),
    .io_y_ae(_2_8_io_y_ae),
    .io_y_sw(_2_8_io_y_sw),
    .io_y_sx(_2_8_io_y_sx),
    .io_y_sr(_2_8_io_y_sr),
    .io_y_pw(_2_8_io_y_pw),
    .io_y_px(_2_8_io_y_px),
    .io_y_pr(_2_8_io_y_pr),
    .io_y_pal(_2_8_io_y_pal),
    .io_y_paa(_2_8_io_y_paa),
    .io_y_eff(_2_8_io_y_eff),
    .io_y_c(_2_8_io_y_c)
  );
  _2_1 _2_9 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130533.4]
    .io_x_ppn(_2_9_io_x_ppn),
    .io_x_u(_2_9_io_x_u),
    .io_x_ae(_2_9_io_x_ae),
    .io_x_sw(_2_9_io_x_sw),
    .io_x_sx(_2_9_io_x_sx),
    .io_x_sr(_2_9_io_x_sr),
    .io_x_pw(_2_9_io_x_pw),
    .io_x_px(_2_9_io_x_px),
    .io_x_pr(_2_9_io_x_pr),
    .io_x_pal(_2_9_io_x_pal),
    .io_x_paa(_2_9_io_x_paa),
    .io_x_eff(_2_9_io_x_eff),
    .io_x_c(_2_9_io_x_c),
    .io_y_ppn(_2_9_io_y_ppn),
    .io_y_u(_2_9_io_y_u),
    .io_y_ae(_2_9_io_y_ae),
    .io_y_sw(_2_9_io_y_sw),
    .io_y_sx(_2_9_io_y_sx),
    .io_y_sr(_2_9_io_y_sr),
    .io_y_pw(_2_9_io_y_pw),
    .io_y_px(_2_9_io_y_px),
    .io_y_pr(_2_9_io_y_pr),
    .io_y_pal(_2_9_io_y_pal),
    .io_y_paa(_2_9_io_y_paa),
    .io_y_eff(_2_9_io_y_eff),
    .io_y_c(_2_9_io_y_c)
  );
  _2_1 _2_10 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130580.4]
    .io_x_ppn(_2_10_io_x_ppn),
    .io_x_u(_2_10_io_x_u),
    .io_x_ae(_2_10_io_x_ae),
    .io_x_sw(_2_10_io_x_sw),
    .io_x_sx(_2_10_io_x_sx),
    .io_x_sr(_2_10_io_x_sr),
    .io_x_pw(_2_10_io_x_pw),
    .io_x_px(_2_10_io_x_px),
    .io_x_pr(_2_10_io_x_pr),
    .io_x_pal(_2_10_io_x_pal),
    .io_x_paa(_2_10_io_x_paa),
    .io_x_eff(_2_10_io_x_eff),
    .io_x_c(_2_10_io_x_c),
    .io_y_ppn(_2_10_io_y_ppn),
    .io_y_u(_2_10_io_y_u),
    .io_y_ae(_2_10_io_y_ae),
    .io_y_sw(_2_10_io_y_sw),
    .io_y_sx(_2_10_io_y_sx),
    .io_y_sr(_2_10_io_y_sr),
    .io_y_pw(_2_10_io_y_pw),
    .io_y_px(_2_10_io_y_px),
    .io_y_pr(_2_10_io_y_pr),
    .io_y_pal(_2_10_io_y_pal),
    .io_y_paa(_2_10_io_y_paa),
    .io_y_eff(_2_10_io_y_eff),
    .io_y_c(_2_10_io_y_c)
  );
  _2_1 _2_11 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130627.4]
    .io_x_ppn(_2_11_io_x_ppn),
    .io_x_u(_2_11_io_x_u),
    .io_x_ae(_2_11_io_x_ae),
    .io_x_sw(_2_11_io_x_sw),
    .io_x_sx(_2_11_io_x_sx),
    .io_x_sr(_2_11_io_x_sr),
    .io_x_pw(_2_11_io_x_pw),
    .io_x_px(_2_11_io_x_px),
    .io_x_pr(_2_11_io_x_pr),
    .io_x_pal(_2_11_io_x_pal),
    .io_x_paa(_2_11_io_x_paa),
    .io_x_eff(_2_11_io_x_eff),
    .io_x_c(_2_11_io_x_c),
    .io_y_ppn(_2_11_io_y_ppn),
    .io_y_u(_2_11_io_y_u),
    .io_y_ae(_2_11_io_y_ae),
    .io_y_sw(_2_11_io_y_sw),
    .io_y_sx(_2_11_io_y_sx),
    .io_y_sr(_2_11_io_y_sr),
    .io_y_pw(_2_11_io_y_pw),
    .io_y_px(_2_11_io_y_px),
    .io_y_pr(_2_11_io_y_pr),
    .io_y_pal(_2_11_io_y_pal),
    .io_y_paa(_2_11_io_y_paa),
    .io_y_eff(_2_11_io_y_eff),
    .io_y_c(_2_11_io_y_c)
  );
  _2_1 _2_12 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130674.4]
    .io_x_ppn(_2_12_io_x_ppn),
    .io_x_u(_2_12_io_x_u),
    .io_x_ae(_2_12_io_x_ae),
    .io_x_sw(_2_12_io_x_sw),
    .io_x_sx(_2_12_io_x_sx),
    .io_x_sr(_2_12_io_x_sr),
    .io_x_pw(_2_12_io_x_pw),
    .io_x_px(_2_12_io_x_px),
    .io_x_pr(_2_12_io_x_pr),
    .io_x_pal(_2_12_io_x_pal),
    .io_x_paa(_2_12_io_x_paa),
    .io_x_eff(_2_12_io_x_eff),
    .io_x_c(_2_12_io_x_c),
    .io_y_ppn(_2_12_io_y_ppn),
    .io_y_u(_2_12_io_y_u),
    .io_y_ae(_2_12_io_y_ae),
    .io_y_sw(_2_12_io_y_sw),
    .io_y_sx(_2_12_io_y_sx),
    .io_y_sr(_2_12_io_y_sr),
    .io_y_pw(_2_12_io_y_pw),
    .io_y_px(_2_12_io_y_px),
    .io_y_pr(_2_12_io_y_pr),
    .io_y_pal(_2_12_io_y_pal),
    .io_y_paa(_2_12_io_y_paa),
    .io_y_eff(_2_12_io_y_eff),
    .io_y_c(_2_12_io_y_c)
  );
  _2_1 _2_13 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@130721.4]
    .io_x_ppn(_2_13_io_x_ppn),
    .io_x_u(_2_13_io_x_u),
    .io_x_ae(_2_13_io_x_ae),
    .io_x_sw(_2_13_io_x_sw),
    .io_x_sx(_2_13_io_x_sx),
    .io_x_sr(_2_13_io_x_sr),
    .io_x_pw(_2_13_io_x_pw),
    .io_x_px(_2_13_io_x_px),
    .io_x_pr(_2_13_io_x_pr),
    .io_x_pal(_2_13_io_x_pal),
    .io_x_paa(_2_13_io_x_paa),
    .io_x_eff(_2_13_io_x_eff),
    .io_x_c(_2_13_io_x_c),
    .io_y_ppn(_2_13_io_y_ppn),
    .io_y_u(_2_13_io_y_u),
    .io_y_ae(_2_13_io_y_ae),
    .io_y_sw(_2_13_io_y_sw),
    .io_y_sx(_2_13_io_y_sx),
    .io_y_sr(_2_13_io_y_sr),
    .io_y_pw(_2_13_io_y_pw),
    .io_y_px(_2_13_io_y_px),
    .io_y_pr(_2_13_io_y_pr),
    .io_y_pal(_2_13_io_y_pal),
    .io_y_paa(_2_13_io_y_paa),
    .io_y_eff(_2_13_io_y_eff),
    .io_y_c(_2_13_io_y_c)
  );
  _2_1 _2_14 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131186.4]
    .io_x_ppn(_2_14_io_x_ppn),
    .io_x_u(_2_14_io_x_u),
    .io_x_ae(_2_14_io_x_ae),
    .io_x_sw(_2_14_io_x_sw),
    .io_x_sx(_2_14_io_x_sx),
    .io_x_sr(_2_14_io_x_sr),
    .io_x_pw(_2_14_io_x_pw),
    .io_x_px(_2_14_io_x_px),
    .io_x_pr(_2_14_io_x_pr),
    .io_x_pal(_2_14_io_x_pal),
    .io_x_paa(_2_14_io_x_paa),
    .io_x_eff(_2_14_io_x_eff),
    .io_x_c(_2_14_io_x_c),
    .io_y_ppn(_2_14_io_y_ppn),
    .io_y_u(_2_14_io_y_u),
    .io_y_ae(_2_14_io_y_ae),
    .io_y_sw(_2_14_io_y_sw),
    .io_y_sx(_2_14_io_y_sx),
    .io_y_sr(_2_14_io_y_sr),
    .io_y_pw(_2_14_io_y_pw),
    .io_y_px(_2_14_io_y_px),
    .io_y_pr(_2_14_io_y_pr),
    .io_y_pal(_2_14_io_y_pal),
    .io_y_paa(_2_14_io_y_paa),
    .io_y_eff(_2_14_io_y_eff),
    .io_y_c(_2_14_io_y_c)
  );
  _2_1 _2_15 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131227.4]
    .io_x_ppn(_2_15_io_x_ppn),
    .io_x_u(_2_15_io_x_u),
    .io_x_ae(_2_15_io_x_ae),
    .io_x_sw(_2_15_io_x_sw),
    .io_x_sx(_2_15_io_x_sx),
    .io_x_sr(_2_15_io_x_sr),
    .io_x_pw(_2_15_io_x_pw),
    .io_x_px(_2_15_io_x_px),
    .io_x_pr(_2_15_io_x_pr),
    .io_x_pal(_2_15_io_x_pal),
    .io_x_paa(_2_15_io_x_paa),
    .io_x_eff(_2_15_io_x_eff),
    .io_x_c(_2_15_io_x_c),
    .io_y_ppn(_2_15_io_y_ppn),
    .io_y_u(_2_15_io_y_u),
    .io_y_ae(_2_15_io_y_ae),
    .io_y_sw(_2_15_io_y_sw),
    .io_y_sx(_2_15_io_y_sx),
    .io_y_sr(_2_15_io_y_sr),
    .io_y_pw(_2_15_io_y_pw),
    .io_y_px(_2_15_io_y_px),
    .io_y_pr(_2_15_io_y_pr),
    .io_y_pal(_2_15_io_y_pal),
    .io_y_paa(_2_15_io_y_paa),
    .io_y_eff(_2_15_io_y_eff),
    .io_y_c(_2_15_io_y_c)
  );
  _2_1 _2_16 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131268.4]
    .io_x_ppn(_2_16_io_x_ppn),
    .io_x_u(_2_16_io_x_u),
    .io_x_ae(_2_16_io_x_ae),
    .io_x_sw(_2_16_io_x_sw),
    .io_x_sx(_2_16_io_x_sx),
    .io_x_sr(_2_16_io_x_sr),
    .io_x_pw(_2_16_io_x_pw),
    .io_x_px(_2_16_io_x_px),
    .io_x_pr(_2_16_io_x_pr),
    .io_x_pal(_2_16_io_x_pal),
    .io_x_paa(_2_16_io_x_paa),
    .io_x_eff(_2_16_io_x_eff),
    .io_x_c(_2_16_io_x_c),
    .io_y_ppn(_2_16_io_y_ppn),
    .io_y_u(_2_16_io_y_u),
    .io_y_ae(_2_16_io_y_ae),
    .io_y_sw(_2_16_io_y_sw),
    .io_y_sx(_2_16_io_y_sx),
    .io_y_sr(_2_16_io_y_sr),
    .io_y_pw(_2_16_io_y_pw),
    .io_y_px(_2_16_io_y_px),
    .io_y_pr(_2_16_io_y_pr),
    .io_y_pal(_2_16_io_y_pal),
    .io_y_paa(_2_16_io_y_paa),
    .io_y_eff(_2_16_io_y_eff),
    .io_y_c(_2_16_io_y_c)
  );
  _2_1 _2_17 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131309.4]
    .io_x_ppn(_2_17_io_x_ppn),
    .io_x_u(_2_17_io_x_u),
    .io_x_ae(_2_17_io_x_ae),
    .io_x_sw(_2_17_io_x_sw),
    .io_x_sx(_2_17_io_x_sx),
    .io_x_sr(_2_17_io_x_sr),
    .io_x_pw(_2_17_io_x_pw),
    .io_x_px(_2_17_io_x_px),
    .io_x_pr(_2_17_io_x_pr),
    .io_x_pal(_2_17_io_x_pal),
    .io_x_paa(_2_17_io_x_paa),
    .io_x_eff(_2_17_io_x_eff),
    .io_x_c(_2_17_io_x_c),
    .io_y_ppn(_2_17_io_y_ppn),
    .io_y_u(_2_17_io_y_u),
    .io_y_ae(_2_17_io_y_ae),
    .io_y_sw(_2_17_io_y_sw),
    .io_y_sx(_2_17_io_y_sx),
    .io_y_sr(_2_17_io_y_sr),
    .io_y_pw(_2_17_io_y_pw),
    .io_y_px(_2_17_io_y_px),
    .io_y_pr(_2_17_io_y_pr),
    .io_y_pal(_2_17_io_y_pal),
    .io_y_paa(_2_17_io_y_paa),
    .io_y_eff(_2_17_io_y_eff),
    .io_y_c(_2_17_io_y_c)
  );
  _2_1 _2_18 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131350.4]
    .io_x_ppn(_2_18_io_x_ppn),
    .io_x_u(_2_18_io_x_u),
    .io_x_ae(_2_18_io_x_ae),
    .io_x_sw(_2_18_io_x_sw),
    .io_x_sx(_2_18_io_x_sx),
    .io_x_sr(_2_18_io_x_sr),
    .io_x_pw(_2_18_io_x_pw),
    .io_x_px(_2_18_io_x_px),
    .io_x_pr(_2_18_io_x_pr),
    .io_x_pal(_2_18_io_x_pal),
    .io_x_paa(_2_18_io_x_paa),
    .io_x_eff(_2_18_io_x_eff),
    .io_x_c(_2_18_io_x_c),
    .io_y_ppn(_2_18_io_y_ppn),
    .io_y_u(_2_18_io_y_u),
    .io_y_ae(_2_18_io_y_ae),
    .io_y_sw(_2_18_io_y_sw),
    .io_y_sx(_2_18_io_y_sx),
    .io_y_sr(_2_18_io_y_sr),
    .io_y_pw(_2_18_io_y_pw),
    .io_y_px(_2_18_io_y_px),
    .io_y_pr(_2_18_io_y_pr),
    .io_y_pal(_2_18_io_y_pal),
    .io_y_paa(_2_18_io_y_paa),
    .io_y_eff(_2_18_io_y_eff),
    .io_y_c(_2_18_io_y_c)
  );
  _2_1 _2_19 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131391.4]
    .io_x_ppn(_2_19_io_x_ppn),
    .io_x_u(_2_19_io_x_u),
    .io_x_ae(_2_19_io_x_ae),
    .io_x_sw(_2_19_io_x_sw),
    .io_x_sx(_2_19_io_x_sx),
    .io_x_sr(_2_19_io_x_sr),
    .io_x_pw(_2_19_io_x_pw),
    .io_x_px(_2_19_io_x_px),
    .io_x_pr(_2_19_io_x_pr),
    .io_x_pal(_2_19_io_x_pal),
    .io_x_paa(_2_19_io_x_paa),
    .io_x_eff(_2_19_io_x_eff),
    .io_x_c(_2_19_io_x_c),
    .io_y_ppn(_2_19_io_y_ppn),
    .io_y_u(_2_19_io_y_u),
    .io_y_ae(_2_19_io_y_ae),
    .io_y_sw(_2_19_io_y_sw),
    .io_y_sx(_2_19_io_y_sx),
    .io_y_sr(_2_19_io_y_sr),
    .io_y_pw(_2_19_io_y_pw),
    .io_y_px(_2_19_io_y_px),
    .io_y_pr(_2_19_io_y_pr),
    .io_y_pal(_2_19_io_y_pal),
    .io_y_paa(_2_19_io_y_paa),
    .io_y_eff(_2_19_io_y_eff),
    .io_y_c(_2_19_io_y_c)
  );
  _2_1 _2_20 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131432.4]
    .io_x_ppn(_2_20_io_x_ppn),
    .io_x_u(_2_20_io_x_u),
    .io_x_ae(_2_20_io_x_ae),
    .io_x_sw(_2_20_io_x_sw),
    .io_x_sx(_2_20_io_x_sx),
    .io_x_sr(_2_20_io_x_sr),
    .io_x_pw(_2_20_io_x_pw),
    .io_x_px(_2_20_io_x_px),
    .io_x_pr(_2_20_io_x_pr),
    .io_x_pal(_2_20_io_x_pal),
    .io_x_paa(_2_20_io_x_paa),
    .io_x_eff(_2_20_io_x_eff),
    .io_x_c(_2_20_io_x_c),
    .io_y_ppn(_2_20_io_y_ppn),
    .io_y_u(_2_20_io_y_u),
    .io_y_ae(_2_20_io_y_ae),
    .io_y_sw(_2_20_io_y_sw),
    .io_y_sx(_2_20_io_y_sx),
    .io_y_sr(_2_20_io_y_sr),
    .io_y_pw(_2_20_io_y_pw),
    .io_y_px(_2_20_io_y_px),
    .io_y_pr(_2_20_io_y_pr),
    .io_y_pal(_2_20_io_y_pal),
    .io_y_paa(_2_20_io_y_paa),
    .io_y_eff(_2_20_io_y_eff),
    .io_y_c(_2_20_io_y_c)
  );
  _2_1 _2_21 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131473.4]
    .io_x_ppn(_2_21_io_x_ppn),
    .io_x_u(_2_21_io_x_u),
    .io_x_ae(_2_21_io_x_ae),
    .io_x_sw(_2_21_io_x_sw),
    .io_x_sx(_2_21_io_x_sx),
    .io_x_sr(_2_21_io_x_sr),
    .io_x_pw(_2_21_io_x_pw),
    .io_x_px(_2_21_io_x_px),
    .io_x_pr(_2_21_io_x_pr),
    .io_x_pal(_2_21_io_x_pal),
    .io_x_paa(_2_21_io_x_paa),
    .io_x_eff(_2_21_io_x_eff),
    .io_x_c(_2_21_io_x_c),
    .io_y_ppn(_2_21_io_y_ppn),
    .io_y_u(_2_21_io_y_u),
    .io_y_ae(_2_21_io_y_ae),
    .io_y_sw(_2_21_io_y_sw),
    .io_y_sx(_2_21_io_y_sx),
    .io_y_sr(_2_21_io_y_sr),
    .io_y_pw(_2_21_io_y_pw),
    .io_y_px(_2_21_io_y_px),
    .io_y_pr(_2_21_io_y_pr),
    .io_y_pal(_2_21_io_y_pal),
    .io_y_paa(_2_21_io_y_paa),
    .io_y_eff(_2_21_io_y_eff),
    .io_y_c(_2_21_io_y_c)
  );
  _2_1 _2_22 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131513.4]
    .io_x_ppn(_2_22_io_x_ppn),
    .io_x_u(_2_22_io_x_u),
    .io_x_ae(_2_22_io_x_ae),
    .io_x_sw(_2_22_io_x_sw),
    .io_x_sx(_2_22_io_x_sx),
    .io_x_sr(_2_22_io_x_sr),
    .io_x_pw(_2_22_io_x_pw),
    .io_x_px(_2_22_io_x_px),
    .io_x_pr(_2_22_io_x_pr),
    .io_x_pal(_2_22_io_x_pal),
    .io_x_paa(_2_22_io_x_paa),
    .io_x_eff(_2_22_io_x_eff),
    .io_x_c(_2_22_io_x_c),
    .io_y_ppn(_2_22_io_y_ppn),
    .io_y_u(_2_22_io_y_u),
    .io_y_ae(_2_22_io_y_ae),
    .io_y_sw(_2_22_io_y_sw),
    .io_y_sx(_2_22_io_y_sx),
    .io_y_sr(_2_22_io_y_sr),
    .io_y_pw(_2_22_io_y_pw),
    .io_y_px(_2_22_io_y_px),
    .io_y_pr(_2_22_io_y_pr),
    .io_y_pal(_2_22_io_y_pal),
    .io_y_paa(_2_22_io_y_paa),
    .io_y_eff(_2_22_io_y_eff),
    .io_y_c(_2_22_io_y_c)
  );
  _2_1 _2_23 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131553.4]
    .io_x_ppn(_2_23_io_x_ppn),
    .io_x_u(_2_23_io_x_u),
    .io_x_ae(_2_23_io_x_ae),
    .io_x_sw(_2_23_io_x_sw),
    .io_x_sx(_2_23_io_x_sx),
    .io_x_sr(_2_23_io_x_sr),
    .io_x_pw(_2_23_io_x_pw),
    .io_x_px(_2_23_io_x_px),
    .io_x_pr(_2_23_io_x_pr),
    .io_x_pal(_2_23_io_x_pal),
    .io_x_paa(_2_23_io_x_paa),
    .io_x_eff(_2_23_io_x_eff),
    .io_x_c(_2_23_io_x_c),
    .io_y_ppn(_2_23_io_y_ppn),
    .io_y_u(_2_23_io_y_u),
    .io_y_ae(_2_23_io_y_ae),
    .io_y_sw(_2_23_io_y_sw),
    .io_y_sx(_2_23_io_y_sx),
    .io_y_sr(_2_23_io_y_sr),
    .io_y_pw(_2_23_io_y_pw),
    .io_y_px(_2_23_io_y_px),
    .io_y_pr(_2_23_io_y_pr),
    .io_y_pal(_2_23_io_y_pal),
    .io_y_paa(_2_23_io_y_paa),
    .io_y_eff(_2_23_io_y_eff),
    .io_y_c(_2_23_io_y_c)
  );
  _2_1 _2_24 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131593.4]
    .io_x_ppn(_2_24_io_x_ppn),
    .io_x_u(_2_24_io_x_u),
    .io_x_ae(_2_24_io_x_ae),
    .io_x_sw(_2_24_io_x_sw),
    .io_x_sx(_2_24_io_x_sx),
    .io_x_sr(_2_24_io_x_sr),
    .io_x_pw(_2_24_io_x_pw),
    .io_x_px(_2_24_io_x_px),
    .io_x_pr(_2_24_io_x_pr),
    .io_x_pal(_2_24_io_x_pal),
    .io_x_paa(_2_24_io_x_paa),
    .io_x_eff(_2_24_io_x_eff),
    .io_x_c(_2_24_io_x_c),
    .io_y_ppn(_2_24_io_y_ppn),
    .io_y_u(_2_24_io_y_u),
    .io_y_ae(_2_24_io_y_ae),
    .io_y_sw(_2_24_io_y_sw),
    .io_y_sx(_2_24_io_y_sx),
    .io_y_sr(_2_24_io_y_sr),
    .io_y_pw(_2_24_io_y_pw),
    .io_y_px(_2_24_io_y_px),
    .io_y_pr(_2_24_io_y_pr),
    .io_y_pal(_2_24_io_y_pal),
    .io_y_paa(_2_24_io_y_paa),
    .io_y_eff(_2_24_io_y_eff),
    .io_y_c(_2_24_io_y_c)
  );
  _2_1 _2_25 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131633.4]
    .io_x_ppn(_2_25_io_x_ppn),
    .io_x_u(_2_25_io_x_u),
    .io_x_ae(_2_25_io_x_ae),
    .io_x_sw(_2_25_io_x_sw),
    .io_x_sx(_2_25_io_x_sx),
    .io_x_sr(_2_25_io_x_sr),
    .io_x_pw(_2_25_io_x_pw),
    .io_x_px(_2_25_io_x_px),
    .io_x_pr(_2_25_io_x_pr),
    .io_x_pal(_2_25_io_x_pal),
    .io_x_paa(_2_25_io_x_paa),
    .io_x_eff(_2_25_io_x_eff),
    .io_x_c(_2_25_io_x_c),
    .io_y_ppn(_2_25_io_y_ppn),
    .io_y_u(_2_25_io_y_u),
    .io_y_ae(_2_25_io_y_ae),
    .io_y_sw(_2_25_io_y_sw),
    .io_y_sx(_2_25_io_y_sx),
    .io_y_sr(_2_25_io_y_sr),
    .io_y_pw(_2_25_io_y_pw),
    .io_y_px(_2_25_io_y_px),
    .io_y_pr(_2_25_io_y_pr),
    .io_y_pal(_2_25_io_y_pal),
    .io_y_paa(_2_25_io_y_paa),
    .io_y_eff(_2_25_io_y_eff),
    .io_y_c(_2_25_io_y_c)
  );
  _2_1 _2_26 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131673.4]
    .io_x_ppn(_2_26_io_x_ppn),
    .io_x_u(_2_26_io_x_u),
    .io_x_ae(_2_26_io_x_ae),
    .io_x_sw(_2_26_io_x_sw),
    .io_x_sx(_2_26_io_x_sx),
    .io_x_sr(_2_26_io_x_sr),
    .io_x_pw(_2_26_io_x_pw),
    .io_x_px(_2_26_io_x_px),
    .io_x_pr(_2_26_io_x_pr),
    .io_x_pal(_2_26_io_x_pal),
    .io_x_paa(_2_26_io_x_paa),
    .io_x_eff(_2_26_io_x_eff),
    .io_x_c(_2_26_io_x_c),
    .io_y_ppn(_2_26_io_y_ppn),
    .io_y_u(_2_26_io_y_u),
    .io_y_ae(_2_26_io_y_ae),
    .io_y_sw(_2_26_io_y_sw),
    .io_y_sx(_2_26_io_y_sx),
    .io_y_sr(_2_26_io_y_sr),
    .io_y_pw(_2_26_io_y_pw),
    .io_y_px(_2_26_io_y_px),
    .io_y_pr(_2_26_io_y_pr),
    .io_y_pal(_2_26_io_y_pal),
    .io_y_paa(_2_26_io_y_paa),
    .io_y_eff(_2_26_io_y_eff),
    .io_y_c(_2_26_io_y_c)
  );
  _2_1 _2_27 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131714.4]
    .io_x_ppn(_2_27_io_x_ppn),
    .io_x_u(_2_27_io_x_u),
    .io_x_ae(_2_27_io_x_ae),
    .io_x_sw(_2_27_io_x_sw),
    .io_x_sx(_2_27_io_x_sx),
    .io_x_sr(_2_27_io_x_sr),
    .io_x_pw(_2_27_io_x_pw),
    .io_x_px(_2_27_io_x_px),
    .io_x_pr(_2_27_io_x_pr),
    .io_x_pal(_2_27_io_x_pal),
    .io_x_paa(_2_27_io_x_paa),
    .io_x_eff(_2_27_io_x_eff),
    .io_x_c(_2_27_io_x_c),
    .io_y_ppn(_2_27_io_y_ppn),
    .io_y_u(_2_27_io_y_u),
    .io_y_ae(_2_27_io_y_ae),
    .io_y_sw(_2_27_io_y_sw),
    .io_y_sx(_2_27_io_y_sx),
    .io_y_sr(_2_27_io_y_sr),
    .io_y_pw(_2_27_io_y_pw),
    .io_y_px(_2_27_io_y_px),
    .io_y_pr(_2_27_io_y_pr),
    .io_y_pal(_2_27_io_y_pal),
    .io_y_paa(_2_27_io_y_paa),
    .io_y_eff(_2_27_io_y_eff),
    .io_y_c(_2_27_io_y_c)
  );
  _2_1 _2_28 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131755.4]
    .io_x_ppn(_2_28_io_x_ppn),
    .io_x_u(_2_28_io_x_u),
    .io_x_ae(_2_28_io_x_ae),
    .io_x_sw(_2_28_io_x_sw),
    .io_x_sx(_2_28_io_x_sx),
    .io_x_sr(_2_28_io_x_sr),
    .io_x_pw(_2_28_io_x_pw),
    .io_x_px(_2_28_io_x_px),
    .io_x_pr(_2_28_io_x_pr),
    .io_x_pal(_2_28_io_x_pal),
    .io_x_paa(_2_28_io_x_paa),
    .io_x_eff(_2_28_io_x_eff),
    .io_x_c(_2_28_io_x_c),
    .io_y_ppn(_2_28_io_y_ppn),
    .io_y_u(_2_28_io_y_u),
    .io_y_ae(_2_28_io_y_ae),
    .io_y_sw(_2_28_io_y_sw),
    .io_y_sx(_2_28_io_y_sx),
    .io_y_sr(_2_28_io_y_sr),
    .io_y_pw(_2_28_io_y_pw),
    .io_y_px(_2_28_io_y_px),
    .io_y_pr(_2_28_io_y_pr),
    .io_y_pal(_2_28_io_y_pal),
    .io_y_paa(_2_28_io_y_paa),
    .io_y_eff(_2_28_io_y_eff),
    .io_y_c(_2_28_io_y_c)
  );
  _2_1 _2_29 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131796.4]
    .io_x_ppn(_2_29_io_x_ppn),
    .io_x_u(_2_29_io_x_u),
    .io_x_ae(_2_29_io_x_ae),
    .io_x_sw(_2_29_io_x_sw),
    .io_x_sx(_2_29_io_x_sx),
    .io_x_sr(_2_29_io_x_sr),
    .io_x_pw(_2_29_io_x_pw),
    .io_x_px(_2_29_io_x_px),
    .io_x_pr(_2_29_io_x_pr),
    .io_x_pal(_2_29_io_x_pal),
    .io_x_paa(_2_29_io_x_paa),
    .io_x_eff(_2_29_io_x_eff),
    .io_x_c(_2_29_io_x_c),
    .io_y_ppn(_2_29_io_y_ppn),
    .io_y_u(_2_29_io_y_u),
    .io_y_ae(_2_29_io_y_ae),
    .io_y_sw(_2_29_io_y_sw),
    .io_y_sx(_2_29_io_y_sx),
    .io_y_sr(_2_29_io_y_sr),
    .io_y_pw(_2_29_io_y_pw),
    .io_y_px(_2_29_io_y_px),
    .io_y_pr(_2_29_io_y_pr),
    .io_y_pal(_2_29_io_y_pal),
    .io_y_paa(_2_29_io_y_paa),
    .io_y_eff(_2_29_io_y_eff),
    .io_y_c(_2_29_io_y_c)
  );
  _2_1 _2_30 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131837.4]
    .io_x_ppn(_2_30_io_x_ppn),
    .io_x_u(_2_30_io_x_u),
    .io_x_ae(_2_30_io_x_ae),
    .io_x_sw(_2_30_io_x_sw),
    .io_x_sx(_2_30_io_x_sx),
    .io_x_sr(_2_30_io_x_sr),
    .io_x_pw(_2_30_io_x_pw),
    .io_x_px(_2_30_io_x_px),
    .io_x_pr(_2_30_io_x_pr),
    .io_x_pal(_2_30_io_x_pal),
    .io_x_paa(_2_30_io_x_paa),
    .io_x_eff(_2_30_io_x_eff),
    .io_x_c(_2_30_io_x_c),
    .io_y_ppn(_2_30_io_y_ppn),
    .io_y_u(_2_30_io_y_u),
    .io_y_ae(_2_30_io_y_ae),
    .io_y_sw(_2_30_io_y_sw),
    .io_y_sx(_2_30_io_y_sx),
    .io_y_sr(_2_30_io_y_sr),
    .io_y_pw(_2_30_io_y_pw),
    .io_y_px(_2_30_io_y_px),
    .io_y_pr(_2_30_io_y_pr),
    .io_y_pal(_2_30_io_y_pal),
    .io_y_paa(_2_30_io_y_paa),
    .io_y_eff(_2_30_io_y_eff),
    .io_y_c(_2_30_io_y_c)
  );
  _2_1 _2_31 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131878.4]
    .io_x_ppn(_2_31_io_x_ppn),
    .io_x_u(_2_31_io_x_u),
    .io_x_ae(_2_31_io_x_ae),
    .io_x_sw(_2_31_io_x_sw),
    .io_x_sx(_2_31_io_x_sx),
    .io_x_sr(_2_31_io_x_sr),
    .io_x_pw(_2_31_io_x_pw),
    .io_x_px(_2_31_io_x_px),
    .io_x_pr(_2_31_io_x_pr),
    .io_x_pal(_2_31_io_x_pal),
    .io_x_paa(_2_31_io_x_paa),
    .io_x_eff(_2_31_io_x_eff),
    .io_x_c(_2_31_io_x_c),
    .io_y_ppn(_2_31_io_y_ppn),
    .io_y_u(_2_31_io_y_u),
    .io_y_ae(_2_31_io_y_ae),
    .io_y_sw(_2_31_io_y_sw),
    .io_y_sx(_2_31_io_y_sx),
    .io_y_sr(_2_31_io_y_sr),
    .io_y_pw(_2_31_io_y_pw),
    .io_y_px(_2_31_io_y_px),
    .io_y_pr(_2_31_io_y_pr),
    .io_y_pal(_2_31_io_y_pal),
    .io_y_paa(_2_31_io_y_paa),
    .io_y_eff(_2_31_io_y_eff),
    .io_y_c(_2_31_io_y_c)
  );
  _2_1 _2_32 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131919.4]
    .io_x_ppn(_2_32_io_x_ppn),
    .io_x_u(_2_32_io_x_u),
    .io_x_ae(_2_32_io_x_ae),
    .io_x_sw(_2_32_io_x_sw),
    .io_x_sx(_2_32_io_x_sx),
    .io_x_sr(_2_32_io_x_sr),
    .io_x_pw(_2_32_io_x_pw),
    .io_x_px(_2_32_io_x_px),
    .io_x_pr(_2_32_io_x_pr),
    .io_x_pal(_2_32_io_x_pal),
    .io_x_paa(_2_32_io_x_paa),
    .io_x_eff(_2_32_io_x_eff),
    .io_x_c(_2_32_io_x_c),
    .io_y_ppn(_2_32_io_y_ppn),
    .io_y_u(_2_32_io_y_u),
    .io_y_ae(_2_32_io_y_ae),
    .io_y_sw(_2_32_io_y_sw),
    .io_y_sx(_2_32_io_y_sx),
    .io_y_sr(_2_32_io_y_sr),
    .io_y_pw(_2_32_io_y_pw),
    .io_y_px(_2_32_io_y_px),
    .io_y_pr(_2_32_io_y_pr),
    .io_y_pal(_2_32_io_y_pal),
    .io_y_paa(_2_32_io_y_paa),
    .io_y_eff(_2_32_io_y_eff),
    .io_y_c(_2_32_io_y_c)
  );
  _2_1 _2_33 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@131960.4]
    .io_x_ppn(_2_33_io_x_ppn),
    .io_x_u(_2_33_io_x_u),
    .io_x_ae(_2_33_io_x_ae),
    .io_x_sw(_2_33_io_x_sw),
    .io_x_sx(_2_33_io_x_sx),
    .io_x_sr(_2_33_io_x_sr),
    .io_x_pw(_2_33_io_x_pw),
    .io_x_px(_2_33_io_x_px),
    .io_x_pr(_2_33_io_x_pr),
    .io_x_pal(_2_33_io_x_pal),
    .io_x_paa(_2_33_io_x_paa),
    .io_x_eff(_2_33_io_x_eff),
    .io_x_c(_2_33_io_x_c),
    .io_y_ppn(_2_33_io_y_ppn),
    .io_y_u(_2_33_io_y_u),
    .io_y_ae(_2_33_io_y_ae),
    .io_y_sw(_2_33_io_y_sw),
    .io_y_sx(_2_33_io_y_sx),
    .io_y_sr(_2_33_io_y_sr),
    .io_y_pw(_2_33_io_y_pw),
    .io_y_px(_2_33_io_y_px),
    .io_y_pr(_2_33_io_y_pr),
    .io_y_pal(_2_33_io_y_pal),
    .io_y_paa(_2_33_io_y_paa),
    .io_y_eff(_2_33_io_y_eff),
    .io_y_c(_2_33_io_y_c)
  );
  _2_1 _2_34 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132001.4]
    .io_x_ppn(_2_34_io_x_ppn),
    .io_x_u(_2_34_io_x_u),
    .io_x_ae(_2_34_io_x_ae),
    .io_x_sw(_2_34_io_x_sw),
    .io_x_sx(_2_34_io_x_sx),
    .io_x_sr(_2_34_io_x_sr),
    .io_x_pw(_2_34_io_x_pw),
    .io_x_px(_2_34_io_x_px),
    .io_x_pr(_2_34_io_x_pr),
    .io_x_pal(_2_34_io_x_pal),
    .io_x_paa(_2_34_io_x_paa),
    .io_x_eff(_2_34_io_x_eff),
    .io_x_c(_2_34_io_x_c),
    .io_y_ppn(_2_34_io_y_ppn),
    .io_y_u(_2_34_io_y_u),
    .io_y_ae(_2_34_io_y_ae),
    .io_y_sw(_2_34_io_y_sw),
    .io_y_sx(_2_34_io_y_sx),
    .io_y_sr(_2_34_io_y_sr),
    .io_y_pw(_2_34_io_y_pw),
    .io_y_px(_2_34_io_y_px),
    .io_y_pr(_2_34_io_y_pr),
    .io_y_pal(_2_34_io_y_pal),
    .io_y_paa(_2_34_io_y_paa),
    .io_y_eff(_2_34_io_y_eff),
    .io_y_c(_2_34_io_y_c)
  );
  _2_1 _2_35 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132041.4]
    .io_x_ppn(_2_35_io_x_ppn),
    .io_x_u(_2_35_io_x_u),
    .io_x_ae(_2_35_io_x_ae),
    .io_x_sw(_2_35_io_x_sw),
    .io_x_sx(_2_35_io_x_sx),
    .io_x_sr(_2_35_io_x_sr),
    .io_x_pw(_2_35_io_x_pw),
    .io_x_px(_2_35_io_x_px),
    .io_x_pr(_2_35_io_x_pr),
    .io_x_pal(_2_35_io_x_pal),
    .io_x_paa(_2_35_io_x_paa),
    .io_x_eff(_2_35_io_x_eff),
    .io_x_c(_2_35_io_x_c),
    .io_y_ppn(_2_35_io_y_ppn),
    .io_y_u(_2_35_io_y_u),
    .io_y_ae(_2_35_io_y_ae),
    .io_y_sw(_2_35_io_y_sw),
    .io_y_sx(_2_35_io_y_sx),
    .io_y_sr(_2_35_io_y_sr),
    .io_y_pw(_2_35_io_y_pw),
    .io_y_px(_2_35_io_y_px),
    .io_y_pr(_2_35_io_y_pr),
    .io_y_pal(_2_35_io_y_pal),
    .io_y_paa(_2_35_io_y_paa),
    .io_y_eff(_2_35_io_y_eff),
    .io_y_c(_2_35_io_y_c)
  );
  _2_1 _2_36 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132081.4]
    .io_x_ppn(_2_36_io_x_ppn),
    .io_x_u(_2_36_io_x_u),
    .io_x_ae(_2_36_io_x_ae),
    .io_x_sw(_2_36_io_x_sw),
    .io_x_sx(_2_36_io_x_sx),
    .io_x_sr(_2_36_io_x_sr),
    .io_x_pw(_2_36_io_x_pw),
    .io_x_px(_2_36_io_x_px),
    .io_x_pr(_2_36_io_x_pr),
    .io_x_pal(_2_36_io_x_pal),
    .io_x_paa(_2_36_io_x_paa),
    .io_x_eff(_2_36_io_x_eff),
    .io_x_c(_2_36_io_x_c),
    .io_y_ppn(_2_36_io_y_ppn),
    .io_y_u(_2_36_io_y_u),
    .io_y_ae(_2_36_io_y_ae),
    .io_y_sw(_2_36_io_y_sw),
    .io_y_sx(_2_36_io_y_sx),
    .io_y_sr(_2_36_io_y_sr),
    .io_y_pw(_2_36_io_y_pw),
    .io_y_px(_2_36_io_y_px),
    .io_y_pr(_2_36_io_y_pr),
    .io_y_pal(_2_36_io_y_pal),
    .io_y_paa(_2_36_io_y_paa),
    .io_y_eff(_2_36_io_y_eff),
    .io_y_c(_2_36_io_y_c)
  );
  _2_1 _2_37 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132121.4]
    .io_x_ppn(_2_37_io_x_ppn),
    .io_x_u(_2_37_io_x_u),
    .io_x_ae(_2_37_io_x_ae),
    .io_x_sw(_2_37_io_x_sw),
    .io_x_sx(_2_37_io_x_sx),
    .io_x_sr(_2_37_io_x_sr),
    .io_x_pw(_2_37_io_x_pw),
    .io_x_px(_2_37_io_x_px),
    .io_x_pr(_2_37_io_x_pr),
    .io_x_pal(_2_37_io_x_pal),
    .io_x_paa(_2_37_io_x_paa),
    .io_x_eff(_2_37_io_x_eff),
    .io_x_c(_2_37_io_x_c),
    .io_y_ppn(_2_37_io_y_ppn),
    .io_y_u(_2_37_io_y_u),
    .io_y_ae(_2_37_io_y_ae),
    .io_y_sw(_2_37_io_y_sw),
    .io_y_sx(_2_37_io_y_sx),
    .io_y_sr(_2_37_io_y_sr),
    .io_y_pw(_2_37_io_y_pw),
    .io_y_px(_2_37_io_y_px),
    .io_y_pr(_2_37_io_y_pr),
    .io_y_pal(_2_37_io_y_pal),
    .io_y_paa(_2_37_io_y_paa),
    .io_y_eff(_2_37_io_y_eff),
    .io_y_c(_2_37_io_y_c)
  );
  _2_1 _2_38 ( // @[package.scala 213:21:freechips.rocketchip.system.DefaultRV32Config.fir@132161.4]
    .io_x_ppn(_2_38_io_x_ppn),
    .io_x_u(_2_38_io_x_u),
    .io_x_ae(_2_38_io_x_ae),
    .io_x_sw(_2_38_io_x_sw),
    .io_x_sx(_2_38_io_x_sx),
    .io_x_sr(_2_38_io_x_sr),
    .io_x_pw(_2_38_io_x_pw),
    .io_x_px(_2_38_io_x_px),
    .io_x_pr(_2_38_io_x_pr),
    .io_x_pal(_2_38_io_x_pal),
    .io_x_paa(_2_38_io_x_paa),
    .io_x_eff(_2_38_io_x_eff),
    .io_x_c(_2_38_io_x_c),
    .io_y_ppn(_2_38_io_y_ppn),
    .io_y_u(_2_38_io_y_u),
    .io_y_ae(_2_38_io_y_ae),
    .io_y_sw(_2_38_io_y_sw),
    .io_y_sx(_2_38_io_y_sx),
    .io_y_sr(_2_38_io_y_sr),
    .io_y_pw(_2_38_io_y_pw),
    .io_y_px(_2_38_io_y_px),
    .io_y_pr(_2_38_io_y_pr),
    .io_y_pal(_2_38_io_y_pal),
    .io_y_paa(_2_38_io_y_paa),
    .io_y_eff(_2_38_io_y_eff),
    .io_y_c(_2_38_io_y_c)
  );
  assign priv_s = io_ptw_status_prv[0]; // @[TLB.scala 176:20:freechips.rocketchip.system.DefaultRV32Config.fir@129471.4]
  assign priv_uses_vm = io_ptw_status_prv <= 2'h1; // @[TLB.scala 177:27:freechips.rocketchip.system.DefaultRV32Config.fir@129472.4]
  assign vm_enabled = io_ptw_ptbr_mode & priv_uses_vm; // @[TLB.scala 178:83:freechips.rocketchip.system.DefaultRV32Config.fir@129475.4]
  assign vpn = io_req_bits_vaddr[31:12]; // @[TLB.scala 181:30:freechips.rocketchip.system.DefaultRV32Config.fir@129478.4]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 182:44:freechips.rocketchip.system.DefaultRV32Config.fir@129479.4]
  assign _T_4 = state == 2'h1; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@129481.4]
  assign _T_5 = state == 2'h3; // @[package.scala 15:47:freechips.rocketchip.system.DefaultRV32Config.fir@129482.4]
  assign invalidate_refill = _T_4 | _T_5; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129483.4]
  assign _T_21 = special_entry_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@129514.4]
  assign _T_24 = _2_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@129525.4]
  assign _T_25 = special_entry_level < 1'h1; // @[TLB.scala 121:30:freechips.rocketchip.system.DefaultRV32Config.fir@129526.4]
  assign _T_27 = _T_25 ? vpn : 20'h0; // @[TLB.scala 122:30:freechips.rocketchip.system.DefaultRV32Config.fir@129528.4]
  assign _T_28 = _T_27 | _2_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@129529.4]
  assign _T_29 = _T_28[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@129530.4]
  assign _T_30 = {_T_24,_T_29}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@129531.4]
  assign _T_31 = io_req_bits_vaddr[31:12]; // @[TLB.scala 186:123:freechips.rocketchip.system.DefaultRV32Config.fir@129532.4]
  assign _T_32 = vm_enabled ? _T_30 : _T_31; // @[TLB.scala 186:20:freechips.rocketchip.system.DefaultRV32Config.fir@129533.4]
  assign mpu_ppn = io_ptw_resp_valid ? refill_ppn : _T_32; // @[TLB.scala 185:20:freechips.rocketchip.system.DefaultRV32Config.fir@129534.4]
  assign _T_33 = io_req_bits_vaddr[11:0]; // @[TLB.scala 187:52:freechips.rocketchip.system.DefaultRV32Config.fir@129535.4]
  assign mpu_physaddr = {mpu_ppn,_T_33}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@129536.4]
  assign _T_36 = {io_ptw_status_debug,io_ptw_status_prv}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@129539.4]
  assign mpu_priv = io_ptw_resp_valid ? 3'h1 : _T_36; // @[TLB.scala 188:27:freechips.rocketchip.system.DefaultRV32Config.fir@129540.4]
  assign _T_37 = mpu_physaddr ^ 32'h3000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129556.4]
  assign _T_38 = {1'b0,$signed(_T_37)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129557.4]
  assign _T_39 = $signed(_T_38) & $signed(-33'sh1000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129558.4]
  assign _T_40 = $signed(_T_39); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129559.4]
  assign _T_41 = $signed(_T_40) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129560.4]
  assign _T_42 = mpu_physaddr ^ 32'hc000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129561.4]
  assign _T_43 = {1'b0,$signed(_T_42)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129562.4]
  assign _T_44 = $signed(_T_43) & $signed(-33'sh4000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129563.4]
  assign _T_45 = $signed(_T_44); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129564.4]
  assign _T_46 = $signed(_T_45) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129565.4]
  assign _T_47 = mpu_physaddr ^ 32'h2000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129566.4]
  assign _T_48 = {1'b0,$signed(_T_47)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129567.4]
  assign _T_49 = $signed(_T_48) & $signed(-33'sh10000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129568.4]
  assign _T_50 = $signed(_T_49); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129569.4]
  assign _T_51 = $signed(_T_50) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129570.4]
  assign _T_53 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129572.4]
  assign _T_54 = $signed(_T_53) & $signed(-33'sh1000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129573.4]
  assign _T_55 = $signed(_T_54); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129574.4]
  assign _T_56 = $signed(_T_55) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129575.4]
  assign _T_57 = mpu_physaddr ^ 32'h10000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129576.4]
  assign _T_58 = {1'b0,$signed(_T_57)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129577.4]
  assign _T_59 = $signed(_T_58) & $signed(-33'sh10000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129578.4]
  assign _T_60 = $signed(_T_59); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129579.4]
  assign _T_61 = $signed(_T_60) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129580.4]
  assign _T_62 = mpu_physaddr ^ 32'h80000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129581.4]
  assign _T_63 = {1'b0,$signed(_T_62)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129582.4]
  assign _T_64 = $signed(_T_63) & $signed(-33'sh10000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129583.4]
  assign _T_65 = $signed(_T_64); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129584.4]
  assign _T_66 = $signed(_T_65) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129585.4]
  assign _T_67 = mpu_physaddr ^ 32'h60000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129586.4]
  assign _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129587.4]
  assign _T_69 = $signed(_T_68) & $signed(-33'sh20000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129588.4]
  assign _T_70 = $signed(_T_69); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129589.4]
  assign _T_71 = $signed(_T_70) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129590.4]
  assign _T_73 = _T_41 | _T_46; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129600.4]
  assign _T_74 = _T_73 | _T_51; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129601.4]
  assign _T_75 = _T_74 | _T_56; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129602.4]
  assign _T_76 = _T_75 | _T_61; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129603.4]
  assign _T_77 = _T_76 | _T_66; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129604.4]
  assign legal_address = _T_77 | _T_71; // @[TLB.scala 194:67:freechips.rocketchip.system.DefaultRV32Config.fir@129605.4]
  assign _T_85 = $signed(_T_63) & $signed(33'sh80000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129613.4]
  assign _T_86 = $signed(_T_85); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129614.4]
  assign _T_87 = $signed(_T_86) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129615.4]
  assign cacheable = legal_address & _T_87; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129621.4]
  assign _T_142 = mpu_physaddr ^ 32'h8000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129673.4]
  assign _T_143 = {1'b0,$signed(_T_142)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129674.4]
  assign _T_144 = $signed(_T_143) & $signed(33'shc8000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129675.4]
  assign _T_145 = $signed(_T_144); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129676.4]
  assign _T_146 = $signed(_T_145) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129677.4]
  assign _T_163 = $signed(_T_53) & $signed(33'shc8010000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129694.4]
  assign _T_164 = $signed(_T_163); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129695.4]
  assign _T_165 = $signed(_T_164) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129696.4]
  assign _T_172 = _T_165 | _T_146; // @[TLBPermissions.scala 82:66:freechips.rocketchip.system.DefaultRV32Config.fir@129703.4]
  assign _T_185 = mpu_priv <= 3'h3; // @[TLB.scala 199:39:freechips.rocketchip.system.DefaultRV32Config.fir@129716.4]
  assign deny_access_to_debug = _T_185 & _T_56; // @[TLB.scala 199:48:freechips.rocketchip.system.DefaultRV32Config.fir@129722.4]
  assign _T_197 = deny_access_to_debug == 1'h0; // @[TLB.scala 200:44:freechips.rocketchip.system.DefaultRV32Config.fir@129729.4]
  assign _T_198 = legal_address & _T_197; // @[TLB.scala 200:41:freechips.rocketchip.system.DefaultRV32Config.fir@129730.4]
  assign prot_r = _T_198 & pmp_io_r; // @[TLB.scala 200:66:freechips.rocketchip.system.DefaultRV32Config.fir@129731.4]
  assign _T_211 = $signed(_T_63) & $signed(33'shc0000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129744.4]
  assign _T_212 = $signed(_T_211); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129745.4]
  assign _T_213 = $signed(_T_212) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129746.4]
  assign _T_214 = mpu_physaddr ^ 32'h40000000; // @[Parameters.scala 125:31:freechips.rocketchip.system.DefaultRV32Config.fir@129747.4]
  assign _T_215 = {1'b0,$signed(_T_214)}; // @[Parameters.scala 125:49:freechips.rocketchip.system.DefaultRV32Config.fir@129748.4]
  assign _T_216 = $signed(_T_215) & $signed(33'shc0000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129749.4]
  assign _T_217 = $signed(_T_216); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129750.4]
  assign _T_218 = $signed(_T_217) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129751.4]
  assign _T_220 = _T_172 | _T_213; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129753.4]
  assign _T_221 = _T_220 | _T_218; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129754.4]
  assign _T_231 = legal_address & _T_221; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129765.4]
  assign _T_233 = _T_231 & _T_197; // @[TLB.scala 201:45:freechips.rocketchip.system.DefaultRV32Config.fir@129767.4]
  assign prot_w = _T_233 & pmp_io_w; // @[TLB.scala 201:70:freechips.rocketchip.system.DefaultRV32Config.fir@129768.4]
  assign prot_al = legal_address & _T_172; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129802.4]
  assign _T_300 = $signed(_T_53) & $signed(33'shca000000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129839.4]
  assign _T_301 = $signed(_T_300); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129840.4]
  assign _T_302 = $signed(_T_301) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129841.4]
  assign _T_313 = _T_302 | _T_213; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129852.4]
  assign _T_314 = _T_313 | _T_218; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129853.4]
  assign _T_330 = legal_address & _T_314; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129870.4]
  assign _T_332 = _T_330 & _T_197; // @[TLB.scala 204:40:freechips.rocketchip.system.DefaultRV32Config.fir@129872.4]
  assign prot_x = _T_332 & pmp_io_x; // @[TLB.scala 204:65:freechips.rocketchip.system.DefaultRV32Config.fir@129873.4]
  assign _T_357 = $signed(_T_48) & $signed(33'shca010000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129898.4]
  assign _T_358 = $signed(_T_357); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129899.4]
  assign _T_359 = $signed(_T_358) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129900.4]
  assign _T_362 = $signed(_T_53) & $signed(33'shca012000); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129903.4]
  assign _T_363 = $signed(_T_362); // @[Parameters.scala 125:52:freechips.rocketchip.system.DefaultRV32Config.fir@129904.4]
  assign _T_364 = $signed(_T_363) == $signed(33'sh0); // @[Parameters.scala 125:67:freechips.rocketchip.system.DefaultRV32Config.fir@129905.4]
  assign _T_370 = _T_146 | _T_359; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129911.4]
  assign _T_371 = _T_370 | _T_364; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129912.4]
  assign _T_372 = _T_371 | _T_218; // @[Parameters.scala 172:89:freechips.rocketchip.system.DefaultRV32Config.fir@129913.4]
  assign prot_eff = legal_address & _T_372; // @[TLB.scala 196:19:freechips.rocketchip.system.DefaultRV32Config.fir@129919.4]
  assign _T_377 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129920.4]
  assign _T_378 = _T_377 | sectored_entries_0_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129921.4]
  assign _T_379 = _T_378 | sectored_entries_0_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129922.4]
  assign _T_380 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129923.4]
  assign _T_381 = _T_380[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129924.4]
  assign _T_382 = _T_381 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129925.4]
  assign sector_hits_0 = _T_379 & _T_382; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129926.4]
  assign _T_383 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129927.4]
  assign _T_384 = _T_383 | sectored_entries_1_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129928.4]
  assign _T_385 = _T_384 | sectored_entries_1_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129929.4]
  assign _T_386 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129930.4]
  assign _T_387 = _T_386[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129931.4]
  assign _T_388 = _T_387 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129932.4]
  assign sector_hits_1 = _T_385 & _T_388; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129933.4]
  assign _T_389 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129934.4]
  assign _T_390 = _T_389 | sectored_entries_2_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129935.4]
  assign _T_391 = _T_390 | sectored_entries_2_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129936.4]
  assign _T_392 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129937.4]
  assign _T_393 = _T_392[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129938.4]
  assign _T_394 = _T_393 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129939.4]
  assign sector_hits_2 = _T_391 & _T_394; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129940.4]
  assign _T_395 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129941.4]
  assign _T_396 = _T_395 | sectored_entries_3_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129942.4]
  assign _T_397 = _T_396 | sectored_entries_3_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129943.4]
  assign _T_398 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129944.4]
  assign _T_399 = _T_398[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129945.4]
  assign _T_400 = _T_399 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129946.4]
  assign sector_hits_3 = _T_397 & _T_400; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129947.4]
  assign _T_401 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129948.4]
  assign _T_402 = _T_401 | sectored_entries_4_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129949.4]
  assign _T_403 = _T_402 | sectored_entries_4_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129950.4]
  assign _T_404 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129951.4]
  assign _T_405 = _T_404[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129952.4]
  assign _T_406 = _T_405 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129953.4]
  assign sector_hits_4 = _T_403 & _T_406; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129954.4]
  assign _T_407 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129955.4]
  assign _T_408 = _T_407 | sectored_entries_5_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129956.4]
  assign _T_409 = _T_408 | sectored_entries_5_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129957.4]
  assign _T_410 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129958.4]
  assign _T_411 = _T_410[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129959.4]
  assign _T_412 = _T_411 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129960.4]
  assign sector_hits_5 = _T_409 & _T_412; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129961.4]
  assign _T_413 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129962.4]
  assign _T_414 = _T_413 | sectored_entries_6_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129963.4]
  assign _T_415 = _T_414 | sectored_entries_6_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129964.4]
  assign _T_416 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129965.4]
  assign _T_417 = _T_416[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129966.4]
  assign _T_418 = _T_417 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129967.4]
  assign sector_hits_6 = _T_415 & _T_418; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129968.4]
  assign _T_419 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129969.4]
  assign _T_420 = _T_419 | sectored_entries_7_valid_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129970.4]
  assign _T_421 = _T_420 | sectored_entries_7_valid_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@129971.4]
  assign _T_422 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 101:43:freechips.rocketchip.system.DefaultRV32Config.fir@129972.4]
  assign _T_423 = _T_422[19:2]; // @[TLB.scala 101:50:freechips.rocketchip.system.DefaultRV32Config.fir@129973.4]
  assign _T_424 = _T_423 == 18'h0; // @[TLB.scala 101:68:freechips.rocketchip.system.DefaultRV32Config.fir@129974.4]
  assign sector_hits_7 = _T_421 & _T_424; // @[TLB.scala 100:42:freechips.rocketchip.system.DefaultRV32Config.fir@129975.4]
  assign _T_427 = superpage_entries_0_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@129978.4]
  assign _T_428 = vpn[19:10]; // @[TLB.scala 108:86:freechips.rocketchip.system.DefaultRV32Config.fir@129979.4]
  assign _T_429 = _T_427 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@129980.4]
  assign superpage_hits_0 = superpage_entries_0_valid_0 & _T_429; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@129982.4]
  assign _T_435 = vpn[9:0]; // @[TLB.scala 108:86:freechips.rocketchip.system.DefaultRV32Config.fir@129986.4]
  assign _T_440 = superpage_entries_1_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@129992.4]
  assign _T_442 = _T_440 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@129994.4]
  assign superpage_hits_1 = superpage_entries_1_valid_0 & _T_442; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@129996.4]
  assign _T_453 = superpage_entries_2_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@130006.4]
  assign _T_455 = _T_453 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@130008.4]
  assign superpage_hits_2 = superpage_entries_2_valid_0 & _T_455; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@130010.4]
  assign _T_466 = superpage_entries_3_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@130020.4]
  assign _T_468 = _T_466 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@130022.4]
  assign superpage_hits_3 = superpage_entries_3_valid_0 & _T_468; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@130024.4]
  assign _T_477 = vpn[1:0]; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@130032.4]
  assign _GEN_1 = 2'h1 == _T_477 ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130036.4]
  assign _GEN_2 = 2'h2 == _T_477 ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130036.4]
  assign _GEN_3 = 2'h3 == _T_477 ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130036.4]
  assign _T_481 = _GEN_3 & _T_382; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130036.4]
  assign hitsVec_0 = vm_enabled & _T_481; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130037.4]
  assign _GEN_5 = 2'h1 == _T_477 ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130042.4]
  assign _GEN_6 = 2'h2 == _T_477 ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130042.4]
  assign _GEN_7 = 2'h3 == _T_477 ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130042.4]
  assign _T_486 = _GEN_7 & _T_388; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130042.4]
  assign hitsVec_1 = vm_enabled & _T_486; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130043.4]
  assign _GEN_9 = 2'h1 == _T_477 ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130048.4]
  assign _GEN_10 = 2'h2 == _T_477 ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130048.4]
  assign _GEN_11 = 2'h3 == _T_477 ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130048.4]
  assign _T_491 = _GEN_11 & _T_394; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130048.4]
  assign hitsVec_2 = vm_enabled & _T_491; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130049.4]
  assign _GEN_13 = 2'h1 == _T_477 ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130054.4]
  assign _GEN_14 = 2'h2 == _T_477 ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130054.4]
  assign _GEN_15 = 2'h3 == _T_477 ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130054.4]
  assign _T_496 = _GEN_15 & _T_400; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130054.4]
  assign hitsVec_3 = vm_enabled & _T_496; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130055.4]
  assign _GEN_17 = 2'h1 == _T_477 ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130060.4]
  assign _GEN_18 = 2'h2 == _T_477 ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130060.4]
  assign _GEN_19 = 2'h3 == _T_477 ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130060.4]
  assign _T_501 = _GEN_19 & _T_406; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130060.4]
  assign hitsVec_4 = vm_enabled & _T_501; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130061.4]
  assign _GEN_21 = 2'h1 == _T_477 ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130066.4]
  assign _GEN_22 = 2'h2 == _T_477 ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130066.4]
  assign _GEN_23 = 2'h3 == _T_477 ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130066.4]
  assign _T_506 = _GEN_23 & _T_412; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130066.4]
  assign hitsVec_5 = vm_enabled & _T_506; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130067.4]
  assign _GEN_25 = 2'h1 == _T_477 ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130072.4]
  assign _GEN_26 = 2'h2 == _T_477 ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130072.4]
  assign _GEN_27 = 2'h3 == _T_477 ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130072.4]
  assign _T_511 = _GEN_27 & _T_418; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130072.4]
  assign hitsVec_6 = vm_enabled & _T_511; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130073.4]
  assign _GEN_29 = 2'h1 == _T_477 ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130078.4]
  assign _GEN_30 = 2'h2 == _T_477 ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130078.4]
  assign _GEN_31 = 2'h3 == _T_477 ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130078.4]
  assign _T_516 = _GEN_31 & _T_424; // @[TLB.scala 113:20:freechips.rocketchip.system.DefaultRV32Config.fir@130078.4]
  assign hitsVec_7 = vm_enabled & _T_516; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130079.4]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130094.4]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130109.4]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130124.4]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130139.4]
  assign _T_575 = special_entry_tag[19:10]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@130142.4]
  assign _T_577 = _T_575 == _T_428; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@130144.4]
  assign _T_579 = special_entry_valid_0 & _T_577; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@130146.4]
  assign _T_582 = special_entry_tag[9:0]; // @[TLB.scala 108:48:freechips.rocketchip.system.DefaultRV32Config.fir@130149.4]
  assign _T_584 = _T_582 == _T_435; // @[TLB.scala 108:79:freechips.rocketchip.system.DefaultRV32Config.fir@130151.4]
  assign _T_585 = _T_25 | _T_584; // @[TLB.scala 108:42:freechips.rocketchip.system.DefaultRV32Config.fir@130152.4]
  assign _T_586 = _T_579 & _T_585; // @[TLB.scala 108:31:freechips.rocketchip.system.DefaultRV32Config.fir@130153.4]
  assign hitsVec_12 = vm_enabled & _T_586; // @[TLB.scala 209:44:freechips.rocketchip.system.DefaultRV32Config.fir@130154.4]
  assign _T_591 = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130159.4]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_591}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130166.4]
  assign _T_598 = vm_enabled == 1'h0; // @[TLB.scala 211:18:freechips.rocketchip.system.DefaultRV32Config.fir@130167.4]
  assign hits = {_T_598,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_591}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130168.4]
  assign _GEN_33 = 2'h1 == _T_477 ? sectored_entries_0_data_1 : sectored_entries_0_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130175.4]
  assign _GEN_34 = 2'h2 == _T_477 ? sectored_entries_0_data_2 : _GEN_33; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130175.4]
  assign _GEN_35 = 2'h3 == _T_477 ? sectored_entries_0_data_3 : _GEN_34; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130175.4]
  assign _GEN_37 = 2'h1 == _T_477 ? sectored_entries_1_data_1 : sectored_entries_1_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130216.4]
  assign _GEN_38 = 2'h2 == _T_477 ? sectored_entries_1_data_2 : _GEN_37; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130216.4]
  assign _GEN_39 = 2'h3 == _T_477 ? sectored_entries_1_data_3 : _GEN_38; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130216.4]
  assign _GEN_41 = 2'h1 == _T_477 ? sectored_entries_2_data_1 : sectored_entries_2_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130257.4]
  assign _GEN_42 = 2'h2 == _T_477 ? sectored_entries_2_data_2 : _GEN_41; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130257.4]
  assign _GEN_43 = 2'h3 == _T_477 ? sectored_entries_2_data_3 : _GEN_42; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130257.4]
  assign _GEN_45 = 2'h1 == _T_477 ? sectored_entries_3_data_1 : sectored_entries_3_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130298.4]
  assign _GEN_46 = 2'h2 == _T_477 ? sectored_entries_3_data_2 : _GEN_45; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130298.4]
  assign _GEN_47 = 2'h3 == _T_477 ? sectored_entries_3_data_3 : _GEN_46; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130298.4]
  assign _GEN_49 = 2'h1 == _T_477 ? sectored_entries_4_data_1 : sectored_entries_4_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130339.4]
  assign _GEN_50 = 2'h2 == _T_477 ? sectored_entries_4_data_2 : _GEN_49; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130339.4]
  assign _GEN_51 = 2'h3 == _T_477 ? sectored_entries_4_data_3 : _GEN_50; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130339.4]
  assign _GEN_53 = 2'h1 == _T_477 ? sectored_entries_5_data_1 : sectored_entries_5_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130380.4]
  assign _GEN_54 = 2'h2 == _T_477 ? sectored_entries_5_data_2 : _GEN_53; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130380.4]
  assign _GEN_55 = 2'h3 == _T_477 ? sectored_entries_5_data_3 : _GEN_54; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130380.4]
  assign _GEN_57 = 2'h1 == _T_477 ? sectored_entries_6_data_1 : sectored_entries_6_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130421.4]
  assign _GEN_58 = 2'h2 == _T_477 ? sectored_entries_6_data_2 : _GEN_57; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130421.4]
  assign _GEN_59 = 2'h3 == _T_477 ? sectored_entries_6_data_3 : _GEN_58; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130421.4]
  assign _GEN_61 = 2'h1 == _T_477 ? sectored_entries_7_data_1 : sectored_entries_7_data_0; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130462.4]
  assign _GEN_62 = 2'h2 == _T_477 ? sectored_entries_7_data_2 : _GEN_61; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130462.4]
  assign _GEN_63 = 2'h3 == _T_477 ? sectored_entries_7_data_3 : _GEN_62; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@130462.4]
  assign _T_758 = superpage_entries_0_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@130527.4]
  assign _T_761 = _2_9_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130538.4]
  assign _T_765 = vpn | _2_9_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130542.4]
  assign _T_766 = _T_765[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130543.4]
  assign _T_767 = {_T_761,_T_766}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130544.4]
  assign _T_782 = superpage_entries_1_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@130574.4]
  assign _T_785 = _2_10_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130585.4]
  assign _T_789 = vpn | _2_10_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130589.4]
  assign _T_790 = _T_789[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130590.4]
  assign _T_791 = {_T_785,_T_790}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130591.4]
  assign _T_806 = superpage_entries_2_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@130621.4]
  assign _T_809 = _2_11_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130632.4]
  assign _T_813 = vpn | _2_11_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130636.4]
  assign _T_814 = _T_813[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130637.4]
  assign _T_815 = {_T_809,_T_814}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130638.4]
  assign _T_830 = superpage_entries_3_data_0[12]; // @[TLB.scala 99:79:freechips.rocketchip.system.DefaultRV32Config.fir@130668.4]
  assign _T_833 = _2_12_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130679.4]
  assign _T_837 = vpn | _2_12_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130683.4]
  assign _T_838 = _T_837[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130684.4]
  assign _T_839 = {_T_833,_T_838}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130685.4]
  assign _T_857 = _2_13_io_y_ppn[19:10]; // @[TLB.scala 119:28:freechips.rocketchip.system.DefaultRV32Config.fir@130726.4]
  assign _T_861 = _T_27 | _2_13_io_y_ppn; // @[TLB.scala 122:49:freechips.rocketchip.system.DefaultRV32Config.fir@130730.4]
  assign _T_862 = _T_861[9:0]; // @[TLB.scala 122:60:freechips.rocketchip.system.DefaultRV32Config.fir@130731.4]
  assign _T_863 = {_T_857,_T_862}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@130732.4]
  assign _T_865 = hitsVec_0 ? _2_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130734.4]
  assign _T_866 = hitsVec_1 ? _2_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130735.4]
  assign _T_867 = hitsVec_2 ? _2_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130736.4]
  assign _T_868 = hitsVec_3 ? _2_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130737.4]
  assign _T_869 = hitsVec_4 ? _2_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130738.4]
  assign _T_870 = hitsVec_5 ? _2_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130739.4]
  assign _T_871 = hitsVec_6 ? _2_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130740.4]
  assign _T_872 = hitsVec_7 ? _2_8_io_y_ppn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130741.4]
  assign _T_873 = hitsVec_8 ? _T_767 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130742.4]
  assign _T_874 = hitsVec_9 ? _T_791 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130743.4]
  assign _T_875 = hitsVec_10 ? _T_815 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130744.4]
  assign _T_876 = hitsVec_11 ? _T_839 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130745.4]
  assign _T_877 = hitsVec_12 ? _T_863 : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130746.4]
  assign _T_878 = _T_598 ? vpn : 20'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130747.4]
  assign _T_879 = _T_865 | _T_866; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130748.4]
  assign _T_880 = _T_879 | _T_867; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130749.4]
  assign _T_881 = _T_880 | _T_868; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130750.4]
  assign _T_882 = _T_881 | _T_869; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130751.4]
  assign _T_883 = _T_882 | _T_870; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130752.4]
  assign _T_884 = _T_883 | _T_871; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130753.4]
  assign _T_885 = _T_884 | _T_872; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130754.4]
  assign _T_886 = _T_885 | _T_873; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130755.4]
  assign _T_887 = _T_886 | _T_874; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130756.4]
  assign _T_888 = _T_887 | _T_875; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130757.4]
  assign _T_889 = _T_888 | _T_876; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130758.4]
  assign _T_890 = _T_889 | _T_877; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130759.4]
  assign ppn = _T_890 | _T_878; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@130760.4]
  assign _T_892 = invalidate_refill == 1'h0; // @[TLB.scala 215:22:freechips.rocketchip.system.DefaultRV32Config.fir@130763.4]
  assign _T_893 = io_ptw_resp_valid & _T_892; // @[TLB.scala 215:19:freechips.rocketchip.system.DefaultRV32Config.fir@130764.4]
  assign _T_895 = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 221:25:freechips.rocketchip.system.DefaultRV32Config.fir@130771.6]
  assign _T_896 = io_ptw_resp_bits_pte_w == 1'h0; // @[PTW.scala 68:47:freechips.rocketchip.system.DefaultRV32Config.fir@130774.6]
  assign _T_897 = io_ptw_resp_bits_pte_x & _T_896; // @[PTW.scala 68:44:freechips.rocketchip.system.DefaultRV32Config.fir@130775.6]
  assign _T_898 = io_ptw_resp_bits_pte_r | _T_897; // @[PTW.scala 68:38:freechips.rocketchip.system.DefaultRV32Config.fir@130776.6]
  assign _T_899 = io_ptw_resp_bits_pte_v & _T_898; // @[PTW.scala 68:32:freechips.rocketchip.system.DefaultRV32Config.fir@130777.6]
  assign _T_900 = _T_899 & io_ptw_resp_bits_pte_a; // @[PTW.scala 68:52:freechips.rocketchip.system.DefaultRV32Config.fir@130778.6]
  assign _T_901 = _T_900 & io_ptw_resp_bits_pte_r; // @[PTW.scala 72:35:freechips.rocketchip.system.DefaultRV32Config.fir@130779.6]
  assign _T_907 = _T_900 & io_ptw_resp_bits_pte_w; // @[PTW.scala 73:35:freechips.rocketchip.system.DefaultRV32Config.fir@130786.6]
  assign _T_908 = _T_907 & io_ptw_resp_bits_pte_d; // @[PTW.scala 73:40:freechips.rocketchip.system.DefaultRV32Config.fir@130787.6]
  assign _T_914 = _T_900 & io_ptw_resp_bits_pte_x; // @[PTW.scala 74:35:freechips.rocketchip.system.DefaultRV32Config.fir@130794.6]
  assign _T_915 = io_ptw_resp_bits_homogeneous == 1'h0; // @[TLB.scala 234:37:freechips.rocketchip.system.DefaultRV32Config.fir@130803.6]
  assign _T_923 = {prot_x,prot_r,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 136:26:freechips.rocketchip.system.DefaultRV32Config.fir@130815.8]
  assign _T_931 = {refill_ppn,io_ptw_resp_bits_pte_u,_T_895,io_ptw_resp_bits_ae,_T_908,_T_914,_T_901,prot_w,_T_923}; // @[TLB.scala 136:26:freechips.rocketchip.system.DefaultRV32Config.fir@130823.8]
  assign _T_932 = io_ptw_resp_bits_level < 1'h1; // @[TLB.scala 236:40:freechips.rocketchip.system.DefaultRV32Config.fir@130827.8]
  assign _T_933 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@130829.10]
  assign _GEN_66 = _T_933 | superpage_entries_0_valid_0; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@130830.10]
  assign _T_948 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@130850.10]
  assign _GEN_70 = _T_948 | superpage_entries_1_valid_0; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@130851.10]
  assign _T_963 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@130871.10]
  assign _GEN_74 = _T_963 | superpage_entries_2_valid_0; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@130872.10]
  assign _T_978 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 237:82:freechips.rocketchip.system.DefaultRV32Config.fir@130892.10]
  assign _GEN_78 = _T_978 | superpage_entries_3_valid_0; // @[TLB.scala 237:89:freechips.rocketchip.system.DefaultRV32Config.fir@130893.10]
  assign _T_993 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 241:22:freechips.rocketchip.system.DefaultRV32Config.fir@130915.10]
  assign _T_994 = _T_993 == 3'h0; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@130916.10]
  assign _T_995 = r_sectored_hit == 1'h0; // @[TLB.scala 243:15:freechips.rocketchip.system.DefaultRV32Config.fir@130918.12]
  assign _GEN_80 = _T_995 ? 1'h0 : sectored_entries_0_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130919.12]
  assign _GEN_81 = _T_995 ? 1'h0 : sectored_entries_0_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130919.12]
  assign _GEN_82 = _T_995 ? 1'h0 : sectored_entries_0_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130919.12]
  assign _GEN_83 = _T_995 ? 1'h0 : sectored_entries_0_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130919.12]
  assign _T_996 = r_refill_tag[1:0]; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@130927.12]
  assign _GEN_950 = 2'h0 == _T_996; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  assign _GEN_84 = _GEN_950 | _GEN_80; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  assign _GEN_951 = 2'h1 == _T_996; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  assign _GEN_85 = _GEN_951 | _GEN_81; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  assign _GEN_952 = 2'h2 == _T_996; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  assign _GEN_86 = _GEN_952 | _GEN_82; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  assign _GEN_953 = 2'h3 == _T_996; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  assign _GEN_87 = _GEN_953 | _GEN_83; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130928.12]
  assign _GEN_92 = _T_994 ? _GEN_84 : sectored_entries_0_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130917.10]
  assign _GEN_93 = _T_994 ? _GEN_85 : sectored_entries_0_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130917.10]
  assign _GEN_94 = _T_994 ? _GEN_86 : sectored_entries_0_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130917.10]
  assign _GEN_95 = _T_994 ? _GEN_87 : sectored_entries_0_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130917.10]
  assign _T_1011 = _T_993 == 3'h1; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@130945.10]
  assign _GEN_102 = _T_995 ? 1'h0 : sectored_entries_1_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130948.12]
  assign _GEN_103 = _T_995 ? 1'h0 : sectored_entries_1_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130948.12]
  assign _GEN_104 = _T_995 ? 1'h0 : sectored_entries_1_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130948.12]
  assign _GEN_105 = _T_995 ? 1'h0 : sectored_entries_1_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130948.12]
  assign _GEN_106 = _GEN_950 | _GEN_102; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130957.12]
  assign _GEN_107 = _GEN_951 | _GEN_103; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130957.12]
  assign _GEN_108 = _GEN_952 | _GEN_104; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130957.12]
  assign _GEN_109 = _GEN_953 | _GEN_105; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130957.12]
  assign _GEN_114 = _T_1011 ? _GEN_106 : sectored_entries_1_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130946.10]
  assign _GEN_115 = _T_1011 ? _GEN_107 : sectored_entries_1_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130946.10]
  assign _GEN_116 = _T_1011 ? _GEN_108 : sectored_entries_1_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130946.10]
  assign _GEN_117 = _T_1011 ? _GEN_109 : sectored_entries_1_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130946.10]
  assign _T_1028 = _T_993 == 3'h2; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@130974.10]
  assign _GEN_124 = _T_995 ? 1'h0 : sectored_entries_2_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130977.12]
  assign _GEN_125 = _T_995 ? 1'h0 : sectored_entries_2_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130977.12]
  assign _GEN_126 = _T_995 ? 1'h0 : sectored_entries_2_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130977.12]
  assign _GEN_127 = _T_995 ? 1'h0 : sectored_entries_2_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@130977.12]
  assign _GEN_128 = _GEN_950 | _GEN_124; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130986.12]
  assign _GEN_129 = _GEN_951 | _GEN_125; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130986.12]
  assign _GEN_130 = _GEN_952 | _GEN_126; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130986.12]
  assign _GEN_131 = _GEN_953 | _GEN_127; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@130986.12]
  assign _GEN_136 = _T_1028 ? _GEN_128 : sectored_entries_2_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130975.10]
  assign _GEN_137 = _T_1028 ? _GEN_129 : sectored_entries_2_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130975.10]
  assign _GEN_138 = _T_1028 ? _GEN_130 : sectored_entries_2_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130975.10]
  assign _GEN_139 = _T_1028 ? _GEN_131 : sectored_entries_2_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@130975.10]
  assign _T_1045 = _T_993 == 3'h3; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131003.10]
  assign _GEN_146 = _T_995 ? 1'h0 : sectored_entries_3_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131006.12]
  assign _GEN_147 = _T_995 ? 1'h0 : sectored_entries_3_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131006.12]
  assign _GEN_148 = _T_995 ? 1'h0 : sectored_entries_3_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131006.12]
  assign _GEN_149 = _T_995 ? 1'h0 : sectored_entries_3_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131006.12]
  assign _GEN_150 = _GEN_950 | _GEN_146; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131015.12]
  assign _GEN_151 = _GEN_951 | _GEN_147; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131015.12]
  assign _GEN_152 = _GEN_952 | _GEN_148; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131015.12]
  assign _GEN_153 = _GEN_953 | _GEN_149; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131015.12]
  assign _GEN_158 = _T_1045 ? _GEN_150 : sectored_entries_3_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131004.10]
  assign _GEN_159 = _T_1045 ? _GEN_151 : sectored_entries_3_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131004.10]
  assign _GEN_160 = _T_1045 ? _GEN_152 : sectored_entries_3_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131004.10]
  assign _GEN_161 = _T_1045 ? _GEN_153 : sectored_entries_3_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131004.10]
  assign _T_1062 = _T_993 == 3'h4; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131032.10]
  assign _GEN_168 = _T_995 ? 1'h0 : sectored_entries_4_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131035.12]
  assign _GEN_169 = _T_995 ? 1'h0 : sectored_entries_4_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131035.12]
  assign _GEN_170 = _T_995 ? 1'h0 : sectored_entries_4_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131035.12]
  assign _GEN_171 = _T_995 ? 1'h0 : sectored_entries_4_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131035.12]
  assign _GEN_172 = _GEN_950 | _GEN_168; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131044.12]
  assign _GEN_173 = _GEN_951 | _GEN_169; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131044.12]
  assign _GEN_174 = _GEN_952 | _GEN_170; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131044.12]
  assign _GEN_175 = _GEN_953 | _GEN_171; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131044.12]
  assign _GEN_180 = _T_1062 ? _GEN_172 : sectored_entries_4_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131033.10]
  assign _GEN_181 = _T_1062 ? _GEN_173 : sectored_entries_4_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131033.10]
  assign _GEN_182 = _T_1062 ? _GEN_174 : sectored_entries_4_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131033.10]
  assign _GEN_183 = _T_1062 ? _GEN_175 : sectored_entries_4_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131033.10]
  assign _T_1079 = _T_993 == 3'h5; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131061.10]
  assign _GEN_190 = _T_995 ? 1'h0 : sectored_entries_5_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131064.12]
  assign _GEN_191 = _T_995 ? 1'h0 : sectored_entries_5_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131064.12]
  assign _GEN_192 = _T_995 ? 1'h0 : sectored_entries_5_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131064.12]
  assign _GEN_193 = _T_995 ? 1'h0 : sectored_entries_5_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131064.12]
  assign _GEN_194 = _GEN_950 | _GEN_190; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131073.12]
  assign _GEN_195 = _GEN_951 | _GEN_191; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131073.12]
  assign _GEN_196 = _GEN_952 | _GEN_192; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131073.12]
  assign _GEN_197 = _GEN_953 | _GEN_193; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131073.12]
  assign _GEN_202 = _T_1079 ? _GEN_194 : sectored_entries_5_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131062.10]
  assign _GEN_203 = _T_1079 ? _GEN_195 : sectored_entries_5_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131062.10]
  assign _GEN_204 = _T_1079 ? _GEN_196 : sectored_entries_5_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131062.10]
  assign _GEN_205 = _T_1079 ? _GEN_197 : sectored_entries_5_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131062.10]
  assign _T_1096 = _T_993 == 3'h6; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131090.10]
  assign _GEN_212 = _T_995 ? 1'h0 : sectored_entries_6_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131093.12]
  assign _GEN_213 = _T_995 ? 1'h0 : sectored_entries_6_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131093.12]
  assign _GEN_214 = _T_995 ? 1'h0 : sectored_entries_6_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131093.12]
  assign _GEN_215 = _T_995 ? 1'h0 : sectored_entries_6_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131093.12]
  assign _GEN_216 = _GEN_950 | _GEN_212; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131102.12]
  assign _GEN_217 = _GEN_951 | _GEN_213; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131102.12]
  assign _GEN_218 = _GEN_952 | _GEN_214; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131102.12]
  assign _GEN_219 = _GEN_953 | _GEN_215; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131102.12]
  assign _GEN_224 = _T_1096 ? _GEN_216 : sectored_entries_6_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131091.10]
  assign _GEN_225 = _T_1096 ? _GEN_217 : sectored_entries_6_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131091.10]
  assign _GEN_226 = _T_1096 ? _GEN_218 : sectored_entries_6_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131091.10]
  assign _GEN_227 = _T_1096 ? _GEN_219 : sectored_entries_6_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131091.10]
  assign _T_1113 = _T_993 == 3'h7; // @[TLB.scala 242:65:freechips.rocketchip.system.DefaultRV32Config.fir@131119.10]
  assign _GEN_234 = _T_995 ? 1'h0 : sectored_entries_7_valid_0; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131122.12]
  assign _GEN_235 = _T_995 ? 1'h0 : sectored_entries_7_valid_1; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131122.12]
  assign _GEN_236 = _T_995 ? 1'h0 : sectored_entries_7_valid_2; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131122.12]
  assign _GEN_237 = _T_995 ? 1'h0 : sectored_entries_7_valid_3; // @[TLB.scala 243:32:freechips.rocketchip.system.DefaultRV32Config.fir@131122.12]
  assign _GEN_238 = _GEN_950 | _GEN_234; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131131.12]
  assign _GEN_239 = _GEN_951 | _GEN_235; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131131.12]
  assign _GEN_240 = _GEN_952 | _GEN_236; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131131.12]
  assign _GEN_241 = _GEN_953 | _GEN_237; // @[TLB.scala 135:18:freechips.rocketchip.system.DefaultRV32Config.fir@131131.12]
  assign _GEN_246 = _T_1113 ? _GEN_238 : sectored_entries_7_valid_0; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131120.10]
  assign _GEN_247 = _T_1113 ? _GEN_239 : sectored_entries_7_valid_1; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131120.10]
  assign _GEN_248 = _T_1113 ? _GEN_240 : sectored_entries_7_valid_2; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131120.10]
  assign _GEN_249 = _T_1113 ? _GEN_241 : sectored_entries_7_valid_3; // @[TLB.scala 242:72:freechips.rocketchip.system.DefaultRV32Config.fir@131120.10]
  assign _GEN_258 = _T_932 ? _GEN_66 : superpage_entries_0_valid_0; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_262 = _T_932 ? _GEN_70 : superpage_entries_1_valid_0; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_266 = _T_932 ? _GEN_74 : superpage_entries_2_valid_0; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_270 = _T_932 ? _GEN_78 : superpage_entries_3_valid_0; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_272 = _T_932 ? sectored_entries_0_valid_0 : _GEN_92; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_273 = _T_932 ? sectored_entries_0_valid_1 : _GEN_93; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_274 = _T_932 ? sectored_entries_0_valid_2 : _GEN_94; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_275 = _T_932 ? sectored_entries_0_valid_3 : _GEN_95; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_282 = _T_932 ? sectored_entries_1_valid_0 : _GEN_114; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_283 = _T_932 ? sectored_entries_1_valid_1 : _GEN_115; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_284 = _T_932 ? sectored_entries_1_valid_2 : _GEN_116; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_285 = _T_932 ? sectored_entries_1_valid_3 : _GEN_117; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_292 = _T_932 ? sectored_entries_2_valid_0 : _GEN_136; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_293 = _T_932 ? sectored_entries_2_valid_1 : _GEN_137; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_294 = _T_932 ? sectored_entries_2_valid_2 : _GEN_138; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_295 = _T_932 ? sectored_entries_2_valid_3 : _GEN_139; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_302 = _T_932 ? sectored_entries_3_valid_0 : _GEN_158; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_303 = _T_932 ? sectored_entries_3_valid_1 : _GEN_159; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_304 = _T_932 ? sectored_entries_3_valid_2 : _GEN_160; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_305 = _T_932 ? sectored_entries_3_valid_3 : _GEN_161; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_312 = _T_932 ? sectored_entries_4_valid_0 : _GEN_180; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_313 = _T_932 ? sectored_entries_4_valid_1 : _GEN_181; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_314 = _T_932 ? sectored_entries_4_valid_2 : _GEN_182; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_315 = _T_932 ? sectored_entries_4_valid_3 : _GEN_183; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_322 = _T_932 ? sectored_entries_5_valid_0 : _GEN_202; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_323 = _T_932 ? sectored_entries_5_valid_1 : _GEN_203; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_324 = _T_932 ? sectored_entries_5_valid_2 : _GEN_204; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_325 = _T_932 ? sectored_entries_5_valid_3 : _GEN_205; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_332 = _T_932 ? sectored_entries_6_valid_0 : _GEN_224; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_333 = _T_932 ? sectored_entries_6_valid_1 : _GEN_225; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_334 = _T_932 ? sectored_entries_6_valid_2 : _GEN_226; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_335 = _T_932 ? sectored_entries_6_valid_3 : _GEN_227; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_342 = _T_932 ? sectored_entries_7_valid_0 : _GEN_246; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_343 = _T_932 ? sectored_entries_7_valid_1 : _GEN_247; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_344 = _T_932 ? sectored_entries_7_valid_2 : _GEN_248; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_345 = _T_932 ? sectored_entries_7_valid_3 : _GEN_249; // @[TLB.scala 236:54:freechips.rocketchip.system.DefaultRV32Config.fir@130828.8]
  assign _GEN_354 = _T_915 | special_entry_valid_0; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_358 = _T_915 ? superpage_entries_0_valid_0 : _GEN_258; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_362 = _T_915 ? superpage_entries_1_valid_0 : _GEN_262; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_366 = _T_915 ? superpage_entries_2_valid_0 : _GEN_266; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_370 = _T_915 ? superpage_entries_3_valid_0 : _GEN_270; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_372 = _T_915 ? sectored_entries_0_valid_0 : _GEN_272; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_373 = _T_915 ? sectored_entries_0_valid_1 : _GEN_273; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_374 = _T_915 ? sectored_entries_0_valid_2 : _GEN_274; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_375 = _T_915 ? sectored_entries_0_valid_3 : _GEN_275; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_382 = _T_915 ? sectored_entries_1_valid_0 : _GEN_282; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_383 = _T_915 ? sectored_entries_1_valid_1 : _GEN_283; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_384 = _T_915 ? sectored_entries_1_valid_2 : _GEN_284; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_385 = _T_915 ? sectored_entries_1_valid_3 : _GEN_285; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_392 = _T_915 ? sectored_entries_2_valid_0 : _GEN_292; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_393 = _T_915 ? sectored_entries_2_valid_1 : _GEN_293; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_394 = _T_915 ? sectored_entries_2_valid_2 : _GEN_294; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_395 = _T_915 ? sectored_entries_2_valid_3 : _GEN_295; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_402 = _T_915 ? sectored_entries_3_valid_0 : _GEN_302; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_403 = _T_915 ? sectored_entries_3_valid_1 : _GEN_303; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_404 = _T_915 ? sectored_entries_3_valid_2 : _GEN_304; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_405 = _T_915 ? sectored_entries_3_valid_3 : _GEN_305; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_412 = _T_915 ? sectored_entries_4_valid_0 : _GEN_312; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_413 = _T_915 ? sectored_entries_4_valid_1 : _GEN_313; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_414 = _T_915 ? sectored_entries_4_valid_2 : _GEN_314; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_415 = _T_915 ? sectored_entries_4_valid_3 : _GEN_315; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_422 = _T_915 ? sectored_entries_5_valid_0 : _GEN_322; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_423 = _T_915 ? sectored_entries_5_valid_1 : _GEN_323; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_424 = _T_915 ? sectored_entries_5_valid_2 : _GEN_324; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_425 = _T_915 ? sectored_entries_5_valid_3 : _GEN_325; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_432 = _T_915 ? sectored_entries_6_valid_0 : _GEN_332; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_433 = _T_915 ? sectored_entries_6_valid_1 : _GEN_333; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_434 = _T_915 ? sectored_entries_6_valid_2 : _GEN_334; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_435 = _T_915 ? sectored_entries_6_valid_3 : _GEN_335; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_442 = _T_915 ? sectored_entries_7_valid_0 : _GEN_342; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_443 = _T_915 ? sectored_entries_7_valid_1 : _GEN_343; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_444 = _T_915 ? sectored_entries_7_valid_2 : _GEN_344; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_445 = _T_915 ? sectored_entries_7_valid_3 : _GEN_345; // @[TLB.scala 234:68:freechips.rocketchip.system.DefaultRV32Config.fir@130805.6]
  assign _GEN_454 = _T_893 ? _GEN_354 : special_entry_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_458 = _T_893 ? _GEN_358 : superpage_entries_0_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_462 = _T_893 ? _GEN_362 : superpage_entries_1_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_466 = _T_893 ? _GEN_366 : superpage_entries_2_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_470 = _T_893 ? _GEN_370 : superpage_entries_3_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_472 = _T_893 ? _GEN_372 : sectored_entries_0_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_473 = _T_893 ? _GEN_373 : sectored_entries_0_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_474 = _T_893 ? _GEN_374 : sectored_entries_0_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_475 = _T_893 ? _GEN_375 : sectored_entries_0_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_482 = _T_893 ? _GEN_382 : sectored_entries_1_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_483 = _T_893 ? _GEN_383 : sectored_entries_1_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_484 = _T_893 ? _GEN_384 : sectored_entries_1_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_485 = _T_893 ? _GEN_385 : sectored_entries_1_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_492 = _T_893 ? _GEN_392 : sectored_entries_2_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_493 = _T_893 ? _GEN_393 : sectored_entries_2_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_494 = _T_893 ? _GEN_394 : sectored_entries_2_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_495 = _T_893 ? _GEN_395 : sectored_entries_2_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_502 = _T_893 ? _GEN_402 : sectored_entries_3_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_503 = _T_893 ? _GEN_403 : sectored_entries_3_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_504 = _T_893 ? _GEN_404 : sectored_entries_3_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_505 = _T_893 ? _GEN_405 : sectored_entries_3_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_512 = _T_893 ? _GEN_412 : sectored_entries_4_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_513 = _T_893 ? _GEN_413 : sectored_entries_4_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_514 = _T_893 ? _GEN_414 : sectored_entries_4_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_515 = _T_893 ? _GEN_415 : sectored_entries_4_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_522 = _T_893 ? _GEN_422 : sectored_entries_5_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_523 = _T_893 ? _GEN_423 : sectored_entries_5_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_524 = _T_893 ? _GEN_424 : sectored_entries_5_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_525 = _T_893 ? _GEN_425 : sectored_entries_5_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_532 = _T_893 ? _GEN_432 : sectored_entries_6_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_533 = _T_893 ? _GEN_433 : sectored_entries_6_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_534 = _T_893 ? _GEN_434 : sectored_entries_6_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_535 = _T_893 ? _GEN_435 : sectored_entries_6_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_542 = _T_893 ? _GEN_442 : sectored_entries_7_valid_0; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_543 = _T_893 ? _GEN_443 : sectored_entries_7_valid_1; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_544 = _T_893 ? _GEN_444 : sectored_entries_7_valid_2; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _GEN_545 = _T_893 ? _GEN_445 : sectored_entries_7_valid_3; // @[TLB.scala 215:42:freechips.rocketchip.system.DefaultRV32Config.fir@130765.4]
  assign _T_1575 = {_2_19_io_y_ae,_2_18_io_y_ae,_2_17_io_y_ae,_2_16_io_y_ae,_2_15_io_y_ae,_2_14_io_y_ae}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132170.4]
  assign ptw_ae_array = {1'h0,_2_26_io_y_ae,_2_25_io_y_ae,_2_24_io_y_ae,_2_23_io_y_ae,_2_22_io_y_ae,_2_21_io_y_ae,_2_20_io_y_ae,_T_1575}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132178.4]
  assign _T_1589 = {_2_19_io_y_u,_2_18_io_y_u,_2_17_io_y_u,_2_16_io_y_u,_2_15_io_y_u,_2_14_io_y_u}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132185.4]
  assign _T_1596 = {_2_26_io_y_u,_2_25_io_y_u,_2_24_io_y_u,_2_23_io_y_u,_2_22_io_y_u,_2_21_io_y_u,_2_20_io_y_u,_T_1589}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132192.4]
  assign _T_1610 = ~ _T_1596; // @[TLB.scala 253:98:freechips.rocketchip.system.DefaultRV32Config.fir@132206.4]
  assign priv_x_ok = priv_s ? _T_1610 : _T_1596; // @[TLB.scala 254:22:freechips.rocketchip.system.DefaultRV32Config.fir@132234.4]
  assign _T_1653 = {_2_19_io_y_sx,_2_18_io_y_sx,_2_17_io_y_sx,_2_16_io_y_sx,_2_15_io_y_sx,_2_14_io_y_sx}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132251.4]
  assign _T_1660 = {_2_26_io_y_sx,_2_25_io_y_sx,_2_24_io_y_sx,_2_23_io_y_sx,_2_22_io_y_sx,_2_21_io_y_sx,_2_20_io_y_sx,_T_1653}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132258.4]
  assign _T_1689 = priv_x_ok & _T_1660; // @[TLB.scala 257:39:freechips.rocketchip.system.DefaultRV32Config.fir@132289.4]
  assign x_array = {1'h1,_T_1689}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132290.4]
  assign _T_1704 = ~ ptw_ae_array; // @[TLB.scala 258:89:freechips.rocketchip.system.DefaultRV32Config.fir@132305.4]
  assign _T_1721 = prot_x ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@132324.4]
  assign _T_1726 = {_2_32_io_y_px,_2_31_io_y_px,_2_30_io_y_px,_2_29_io_y_px,_2_28_io_y_px,_2_27_io_y_px}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132329.4]
  assign _T_1733 = {_T_1721,_2_38_io_y_px,_2_37_io_y_px,_2_36_io_y_px,_2_35_io_y_px,_2_34_io_y_px,_2_33_io_y_px,_T_1726}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132336.4]
  assign px_array = _T_1733 & _T_1704; // @[TLB.scala 260:87:freechips.rocketchip.system.DefaultRV32Config.fir@132338.4]
  assign _T_1749 = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@132354.4]
  assign _T_1754 = {_2_32_io_y_c,_2_31_io_y_c,_2_30_io_y_c,_2_29_io_y_c,_2_28_io_y_c,_2_27_io_y_c}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132359.4]
  assign c_array = {_T_1749,_2_38_io_y_c,_2_37_io_y_c,_2_36_io_y_c,_2_35_io_y_c,_2_34_io_y_c,_2_33_io_y_c,_T_1754}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132366.4]
  assign _T_1900 = x_array | ptw_ae_array; // @[TLB.scala 305:33:freechips.rocketchip.system.DefaultRV32Config.fir@132527.4]
  assign pf_inst_array = ~ _T_1900; // @[TLB.scala 305:23:freechips.rocketchip.system.DefaultRV32Config.fir@132528.4]
  assign tlb_hit = real_hits != 13'h0; // @[TLB.scala 307:27:freechips.rocketchip.system.DefaultRV32Config.fir@132529.4]
  assign _T_1903 = tlb_hit == 1'h0; // @[TLB.scala 308:43:freechips.rocketchip.system.DefaultRV32Config.fir@132532.4]
  assign tlb_miss = vm_enabled & _T_1903; // @[TLB.scala 308:40:freechips.rocketchip.system.DefaultRV32Config.fir@132533.4]
  assign _T_1906 = io_req_valid & vm_enabled; // @[TLB.scala 312:22:freechips.rocketchip.system.DefaultRV32Config.fir@132536.4]
  assign _T_1907 = sector_hits_0 | sector_hits_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132538.6]
  assign _T_1908 = _T_1907 | sector_hits_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132539.6]
  assign _T_1909 = _T_1908 | sector_hits_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132540.6]
  assign _T_1910 = _T_1909 | sector_hits_4; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132541.6]
  assign _T_1911 = _T_1910 | sector_hits_5; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132542.6]
  assign _T_1912 = _T_1911 | sector_hits_6; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132543.6]
  assign _T_1913 = _T_1912 | sector_hits_7; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132544.6]
  assign _T_1920 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132552.8]
  assign _T_1921 = _T_1920[7:4]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@132553.8]
  assign _T_1922 = _T_1920[3:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@132554.8]
  assign _T_1923 = _T_1921 != 4'h0; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@132555.8]
  assign _T_1924 = _T_1921 | _T_1922; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@132556.8]
  assign _T_1925 = _T_1924[3:2]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@132557.8]
  assign _T_1926 = _T_1924[1:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@132558.8]
  assign _T_1927 = _T_1925 != 2'h0; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@132559.8]
  assign _T_1928 = _T_1925 | _T_1926; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@132560.8]
  assign _T_1929 = _T_1928[1]; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@132561.8]
  assign _T_1931 = {_T_1923,_T_1927,_T_1929}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132563.8]
  assign _T_1932 = {_T_1904, 1'h0}; // @[Replacement.scala 46:28:freechips.rocketchip.system.DefaultRV32Config.fir@132564.8]
  assign _T_1933 = _T_1931[2]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132565.8]
  assign _T_1934 = _T_1933 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132566.8]
  assign _T_1936 = _T_1932 | 8'h2; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132568.8]
  assign _T_1937 = ~ _T_1932; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132569.8]
  assign _T_1938 = _T_1937 | 8'h2; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132570.8]
  assign _T_1939 = ~ _T_1938; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132571.8]
  assign _T_1940 = _T_1934 ? _T_1936 : _T_1939; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132572.8]
  assign _T_1941 = {1'h1,_T_1933}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132573.8]
  assign _T_1942 = _T_1931[1]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132574.8]
  assign _T_1943 = _T_1942 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132575.8]
  assign _T_1944 = 4'h1 << _T_1941; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132576.8]
  assign _GEN_983 = {{4'd0}, _T_1944}; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132577.8]
  assign _T_1945 = _T_1940 | _GEN_983; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132577.8]
  assign _T_1946 = ~ _T_1940; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132578.8]
  assign _T_1947 = _T_1946 | _GEN_983; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132579.8]
  assign _T_1948 = ~ _T_1947; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132580.8]
  assign _T_1949 = _T_1943 ? _T_1945 : _T_1948; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132581.8]
  assign _T_1950 = {1'h1,_T_1933,_T_1942}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132582.8]
  assign _T_1951 = _T_1931[0]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132583.8]
  assign _T_1952 = _T_1951 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132584.8]
  assign _T_1953 = 8'h1 << _T_1950; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132585.8]
  assign _T_1954 = _T_1949 | _T_1953; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132586.8]
  assign _T_1955 = ~ _T_1949; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132587.8]
  assign _T_1956 = _T_1955 | _T_1953; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132588.8]
  assign _T_1957 = ~ _T_1956; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132589.8]
  assign _T_1958 = _T_1952 ? _T_1954 : _T_1957; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132590.8]
  assign _T_1960 = _T_1958[7:1]; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@132592.8]
  assign _T_1961 = superpage_hits_0 | superpage_hits_1; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132595.6]
  assign _T_1962 = _T_1961 | superpage_hits_2; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132596.6]
  assign _T_1963 = _T_1962 | superpage_hits_3; // @[package.scala 64:59:freechips.rocketchip.system.DefaultRV32Config.fir@132597.6]
  assign _T_1966 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132601.8]
  assign _T_1967 = _T_1966[3:2]; // @[OneHot.scala 30:18:freechips.rocketchip.system.DefaultRV32Config.fir@132602.8]
  assign _T_1968 = _T_1966[1:0]; // @[OneHot.scala 31:18:freechips.rocketchip.system.DefaultRV32Config.fir@132603.8]
  assign _T_1969 = _T_1967 != 2'h0; // @[OneHot.scala 32:14:freechips.rocketchip.system.DefaultRV32Config.fir@132604.8]
  assign _T_1970 = _T_1967 | _T_1968; // @[OneHot.scala 32:28:freechips.rocketchip.system.DefaultRV32Config.fir@132605.8]
  assign _T_1971 = _T_1970[1]; // @[CircuitMath.scala 30:8:freechips.rocketchip.system.DefaultRV32Config.fir@132606.8]
  assign _T_1972 = {_T_1969,_T_1971}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132607.8]
  assign _T_1973 = {_T_1905, 1'h0}; // @[Replacement.scala 46:28:freechips.rocketchip.system.DefaultRV32Config.fir@132608.8]
  assign _T_1974 = _T_1972[1]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132609.8]
  assign _T_1975 = _T_1974 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132610.8]
  assign _T_1977 = _T_1973 | 4'h2; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132612.8]
  assign _T_1978 = ~ _T_1973; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132613.8]
  assign _T_1979 = _T_1978 | 4'h2; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132614.8]
  assign _T_1980 = ~ _T_1979; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132615.8]
  assign _T_1981 = _T_1975 ? _T_1977 : _T_1980; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132616.8]
  assign _T_1982 = {1'h1,_T_1974}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132617.8]
  assign _T_1983 = _T_1972[0]; // @[Replacement.scala 49:20:freechips.rocketchip.system.DefaultRV32Config.fir@132618.8]
  assign _T_1984 = _T_1983 == 1'h0; // @[Replacement.scala 50:43:freechips.rocketchip.system.DefaultRV32Config.fir@132619.8]
  assign _T_1985 = 4'h1 << _T_1982; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132620.8]
  assign _T_1986 = _T_1981 | _T_1985; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132621.8]
  assign _T_1987 = ~ _T_1981; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132622.8]
  assign _T_1988 = _T_1987 | _T_1985; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132623.8]
  assign _T_1989 = ~ _T_1988; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132624.8]
  assign _T_1990 = _T_1984 ? _T_1986 : _T_1989; // @[Replacement.scala 50:37:freechips.rocketchip.system.DefaultRV32Config.fir@132625.8]
  assign _T_1992 = _T_1990[3:1]; // @[package.scala 120:13:freechips.rocketchip.system.DefaultRV32Config.fir@132627.8]
  assign _T_1993 = real_hits[5:0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132631.4]
  assign _T_1994 = _T_1993[2:0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132632.4]
  assign _T_1995 = _T_1994[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132633.4]
  assign _T_1997 = _T_1994[2:1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132635.4]
  assign _T_1998 = _T_1997[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132636.4]
  assign _T_2000 = _T_1997[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132638.4]
  assign _T_2002 = _T_1998 | _T_2000; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132640.4]
  assign _T_2004 = _T_1998 & _T_2000; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132642.4]
  assign _T_2006 = _T_1995 | _T_2002; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132644.4]
  assign _T_2008 = _T_1995 & _T_2002; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132646.4]
  assign _T_2009 = _T_2004 | _T_2008; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132647.4]
  assign _T_2010 = _T_1993[5:3]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132648.4]
  assign _T_2011 = _T_2010[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132649.4]
  assign _T_2013 = _T_2010[2:1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132651.4]
  assign _T_2014 = _T_2013[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132652.4]
  assign _T_2016 = _T_2013[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132654.4]
  assign _T_2018 = _T_2014 | _T_2016; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132656.4]
  assign _T_2020 = _T_2014 & _T_2016; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132658.4]
  assign _T_2022 = _T_2011 | _T_2018; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132660.4]
  assign _T_2024 = _T_2011 & _T_2018; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132662.4]
  assign _T_2025 = _T_2020 | _T_2024; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132663.4]
  assign _T_2026 = _T_2006 | _T_2022; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132664.4]
  assign _T_2027 = _T_2009 | _T_2025; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@132665.4]
  assign _T_2028 = _T_2006 & _T_2022; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132666.4]
  assign _T_2029 = _T_2027 | _T_2028; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132667.4]
  assign _T_2030 = real_hits[12:6]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132668.4]
  assign _T_2031 = _T_2030[2:0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132669.4]
  assign _T_2032 = _T_2031[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132670.4]
  assign _T_2034 = _T_2031[2:1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132672.4]
  assign _T_2035 = _T_2034[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132673.4]
  assign _T_2037 = _T_2034[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132675.4]
  assign _T_2039 = _T_2035 | _T_2037; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132677.4]
  assign _T_2041 = _T_2035 & _T_2037; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132679.4]
  assign _T_2043 = _T_2032 | _T_2039; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132681.4]
  assign _T_2045 = _T_2032 & _T_2039; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132683.4]
  assign _T_2046 = _T_2041 | _T_2045; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132684.4]
  assign _T_2047 = _T_2030[6:3]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132685.4]
  assign _T_2048 = _T_2047[1:0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132686.4]
  assign _T_2049 = _T_2048[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132687.4]
  assign _T_2051 = _T_2048[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132689.4]
  assign _T_2053 = _T_2049 | _T_2051; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132691.4]
  assign _T_2055 = _T_2049 & _T_2051; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132693.4]
  assign _T_2057 = _T_2047[3:2]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132695.4]
  assign _T_2058 = _T_2057[0]; // @[Misc.scala 179:37:freechips.rocketchip.system.DefaultRV32Config.fir@132696.4]
  assign _T_2060 = _T_2057[1]; // @[Misc.scala 180:39:freechips.rocketchip.system.DefaultRV32Config.fir@132698.4]
  assign _T_2062 = _T_2058 | _T_2060; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132700.4]
  assign _T_2064 = _T_2058 & _T_2060; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132702.4]
  assign _T_2066 = _T_2053 | _T_2062; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132704.4]
  assign _T_2067 = _T_2055 | _T_2064; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@132705.4]
  assign _T_2068 = _T_2053 & _T_2062; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132706.4]
  assign _T_2069 = _T_2067 | _T_2068; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132707.4]
  assign _T_2070 = _T_2043 | _T_2066; // @[Misc.scala 181:16:freechips.rocketchip.system.DefaultRV32Config.fir@132708.4]
  assign _T_2071 = _T_2046 | _T_2069; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@132709.4]
  assign _T_2072 = _T_2043 & _T_2066; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132710.4]
  assign _T_2073 = _T_2071 | _T_2072; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132711.4]
  assign _T_2075 = _T_2029 | _T_2073; // @[Misc.scala 181:37:freechips.rocketchip.system.DefaultRV32Config.fir@132713.4]
  assign _T_2076 = _T_2026 & _T_2070; // @[Misc.scala 181:61:freechips.rocketchip.system.DefaultRV32Config.fir@132714.4]
  assign multipleHits = _T_2075 | _T_2076; // @[Misc.scala 181:49:freechips.rocketchip.system.DefaultRV32Config.fir@132715.4]
  assign _T_2086 = pf_inst_array & hits; // @[TLB.scala 327:47:freechips.rocketchip.system.DefaultRV32Config.fir@132728.4]
  assign _T_2093 = ~ px_array; // @[TLB.scala 330:23:freechips.rocketchip.system.DefaultRV32Config.fir@132738.4]
  assign _T_2094 = _T_2093 & hits; // @[TLB.scala 330:33:freechips.rocketchip.system.DefaultRV32Config.fir@132739.4]
  assign _T_2100 = c_array & hits; // @[TLB.scala 334:33:freechips.rocketchip.system.DefaultRV32Config.fir@132749.4]
  assign _T_2107 = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 337:29:freechips.rocketchip.system.DefaultRV32Config.fir@132759.4]
  assign _T_2113 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@132770.4]
  assign _T_2114 = _T_2113 & tlb_miss; // @[TLB.scala 346:25:freechips.rocketchip.system.DefaultRV32Config.fir@132771.4]
  assign _GEN_985 = _T_1973[3:1]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132779.6]
  assign _T_2119 = {{1'd0}, _GEN_985}; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132779.6]
  assign _T_2120 = _T_2119[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132780.6]
  assign _T_2122 = {1'h1,_T_2120}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132782.6]
  assign _T_2126 = _T_1973 >> _T_2122; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132786.6]
  assign _T_2127 = _T_2126[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132787.6]
  assign _T_2129 = {1'h1,_T_2120,_T_2127}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132789.6]
  assign _T_2130 = _T_2129[1:0]; // @[Replacement.scala 63:8:freechips.rocketchip.system.DefaultRV32Config.fir@132790.6]
  assign _T_2133 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132793.6]
  assign _T_2134 = _T_2133 == 4'hf; // @[TLB.scala 394:16:freechips.rocketchip.system.DefaultRV32Config.fir@132794.6]
  assign _T_2135 = ~ _T_2133; // @[TLB.scala 394:43:freechips.rocketchip.system.DefaultRV32Config.fir@132795.6]
  assign _T_2136 = _T_2135[0]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132796.6]
  assign _T_2137 = _T_2135[1]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132797.6]
  assign _T_2138 = _T_2135[2]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132798.6]
  assign _GEN_986 = _T_1932[7:1]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132809.6]
  assign _T_2148 = {{1'd0}, _GEN_986}; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132809.6]
  assign _T_2149 = _T_2148[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132810.6]
  assign _T_2151 = {1'h1,_T_2149}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132812.6]
  assign _T_2155 = _T_1932 >> _T_2151; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132816.6]
  assign _T_2156 = _T_2155[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132817.6]
  assign _T_2158 = {1'h1,_T_2149,_T_2156}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132819.6]
  assign _T_2162 = _T_1932 >> _T_2158; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132823.6]
  assign _T_2163 = _T_2162[0]; // @[Replacement.scala 61:48:freechips.rocketchip.system.DefaultRV32Config.fir@132824.6]
  assign _T_2165 = {1'h1,_T_2149,_T_2156,_T_2163}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132826.6]
  assign _T_2166 = _T_2165[2:0]; // @[Replacement.scala 63:8:freechips.rocketchip.system.DefaultRV32Config.fir@132827.6]
  assign _T_2197 = {_T_421,_T_415,_T_409,_T_403,_T_397,_T_391,_T_385,_T_379}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@132858.6]
  assign _T_2198 = _T_2197 == 8'hff; // @[TLB.scala 394:16:freechips.rocketchip.system.DefaultRV32Config.fir@132859.6]
  assign _T_2199 = ~ _T_2197; // @[TLB.scala 394:43:freechips.rocketchip.system.DefaultRV32Config.fir@132860.6]
  assign _T_2200 = _T_2199[0]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132861.6]
  assign _T_2201 = _T_2199[1]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132862.6]
  assign _T_2202 = _T_2199[2]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132863.6]
  assign _T_2203 = _T_2199[3]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132864.6]
  assign _T_2204 = _T_2199[4]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132865.6]
  assign _T_2205 = _T_2199[5]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132866.6]
  assign _T_2206 = _T_2199[6]; // @[OneHot.scala 47:40:freechips.rocketchip.system.DefaultRV32Config.fir@132867.6]
  assign _T_2243 = state == 2'h2; // @[TLB.scala 360:17:freechips.rocketchip.system.DefaultRV32Config.fir@132919.4]
  assign _T_2244 = _T_2243 & io_sfence_valid; // @[TLB.scala 360:28:freechips.rocketchip.system.DefaultRV32Config.fir@132920.4]
  assign _T_2245 = io_sfence_bits_rs1 == 1'h0; // @[TLB.scala 368:14:freechips.rocketchip.system.DefaultRV32Config.fir@132928.6]
  assign _T_2246 = io_sfence_bits_addr[31:12]; // @[TLB.scala 368:58:freechips.rocketchip.system.DefaultRV32Config.fir@132929.6]
  assign _T_2247 = _T_2246 == vpn; // @[TLB.scala 368:72:freechips.rocketchip.system.DefaultRV32Config.fir@132930.6]
  assign _T_2248 = _T_2245 | _T_2247; // @[TLB.scala 368:34:freechips.rocketchip.system.DefaultRV32Config.fir@132931.6]
  assign _T_2250 = _T_2248 | reset; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@132933.6]
  assign _T_2251 = _T_2250 == 1'h0; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@132934.6]
  assign _T_2257 = _T_380[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@132948.8]
  assign _T_2258 = _T_2257 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@132949.8]
  assign _T_2261 = sectored_entries_0_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@132956.10]
  assign _T_2273 = sectored_entries_0_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@132980.10]
  assign _T_2278 = sectored_entries_0_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@132991.10]
  assign _T_2290 = sectored_entries_0_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133015.10]
  assign _T_2295 = sectored_entries_0_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133026.10]
  assign _T_2307 = sectored_entries_0_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133050.10]
  assign _T_2312 = sectored_entries_0_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133061.10]
  assign _T_2324 = sectored_entries_0_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133085.10]
  assign _T_2395 = _T_2273 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133247.10]
  assign _GEN_648 = _T_2395 ? 1'h0 : _GEN_472; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133248.10]
  assign _T_2396 = _T_2290 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133251.10]
  assign _GEN_649 = _T_2396 ? 1'h0 : _GEN_473; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133252.10]
  assign _T_2397 = _T_2307 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133255.10]
  assign _GEN_650 = _T_2397 ? 1'h0 : _GEN_474; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133256.10]
  assign _T_2398 = _T_2324 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133259.10]
  assign _GEN_651 = _T_2398 ? 1'h0 : _GEN_475; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133260.10]
  assign _GEN_652 = io_sfence_bits_rs2 & _GEN_648; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133106.8]
  assign _GEN_653 = io_sfence_bits_rs2 & _GEN_649; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133106.8]
  assign _GEN_654 = io_sfence_bits_rs2 & _GEN_650; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133106.8]
  assign _GEN_655 = io_sfence_bits_rs2 & _GEN_651; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133106.8]
  assign _T_2404 = _T_386[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@133279.8]
  assign _T_2405 = _T_2404 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@133280.8]
  assign _T_2408 = sectored_entries_1_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133287.10]
  assign _T_2420 = sectored_entries_1_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133311.10]
  assign _T_2425 = sectored_entries_1_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133322.10]
  assign _T_2437 = sectored_entries_1_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133346.10]
  assign _T_2442 = sectored_entries_1_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133357.10]
  assign _T_2454 = sectored_entries_1_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133381.10]
  assign _T_2459 = sectored_entries_1_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133392.10]
  assign _T_2471 = sectored_entries_1_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133416.10]
  assign _T_2542 = _T_2420 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133578.10]
  assign _GEN_676 = _T_2542 ? 1'h0 : _GEN_482; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133579.10]
  assign _T_2543 = _T_2437 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133582.10]
  assign _GEN_677 = _T_2543 ? 1'h0 : _GEN_483; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133583.10]
  assign _T_2544 = _T_2454 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133586.10]
  assign _GEN_678 = _T_2544 ? 1'h0 : _GEN_484; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133587.10]
  assign _T_2545 = _T_2471 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133590.10]
  assign _GEN_679 = _T_2545 ? 1'h0 : _GEN_485; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133591.10]
  assign _GEN_680 = io_sfence_bits_rs2 & _GEN_676; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133437.8]
  assign _GEN_681 = io_sfence_bits_rs2 & _GEN_677; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133437.8]
  assign _GEN_682 = io_sfence_bits_rs2 & _GEN_678; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133437.8]
  assign _GEN_683 = io_sfence_bits_rs2 & _GEN_679; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133437.8]
  assign _T_2551 = _T_392[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@133610.8]
  assign _T_2552 = _T_2551 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@133611.8]
  assign _T_2555 = sectored_entries_2_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133618.10]
  assign _T_2567 = sectored_entries_2_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133642.10]
  assign _T_2572 = sectored_entries_2_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133653.10]
  assign _T_2584 = sectored_entries_2_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133677.10]
  assign _T_2589 = sectored_entries_2_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133688.10]
  assign _T_2601 = sectored_entries_2_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133712.10]
  assign _T_2606 = sectored_entries_2_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133723.10]
  assign _T_2618 = sectored_entries_2_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133747.10]
  assign _T_2689 = _T_2567 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133909.10]
  assign _GEN_704 = _T_2689 ? 1'h0 : _GEN_492; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133910.10]
  assign _T_2690 = _T_2584 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133913.10]
  assign _GEN_705 = _T_2690 ? 1'h0 : _GEN_493; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133914.10]
  assign _T_2691 = _T_2601 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133917.10]
  assign _GEN_706 = _T_2691 ? 1'h0 : _GEN_494; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133918.10]
  assign _T_2692 = _T_2618 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@133921.10]
  assign _GEN_707 = _T_2692 ? 1'h0 : _GEN_495; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@133922.10]
  assign _GEN_708 = io_sfence_bits_rs2 & _GEN_704; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133768.8]
  assign _GEN_709 = io_sfence_bits_rs2 & _GEN_705; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133768.8]
  assign _GEN_710 = io_sfence_bits_rs2 & _GEN_706; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133768.8]
  assign _GEN_711 = io_sfence_bits_rs2 & _GEN_707; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@133768.8]
  assign _T_2698 = _T_398[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@133941.8]
  assign _T_2699 = _T_2698 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@133942.8]
  assign _T_2702 = sectored_entries_3_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133949.10]
  assign _T_2714 = sectored_entries_3_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133973.10]
  assign _T_2719 = sectored_entries_3_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@133984.10]
  assign _T_2731 = sectored_entries_3_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134008.10]
  assign _T_2736 = sectored_entries_3_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134019.10]
  assign _T_2748 = sectored_entries_3_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134043.10]
  assign _T_2753 = sectored_entries_3_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134054.10]
  assign _T_2765 = sectored_entries_3_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134078.10]
  assign _T_2836 = _T_2714 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134240.10]
  assign _GEN_732 = _T_2836 ? 1'h0 : _GEN_502; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134241.10]
  assign _T_2837 = _T_2731 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134244.10]
  assign _GEN_733 = _T_2837 ? 1'h0 : _GEN_503; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134245.10]
  assign _T_2838 = _T_2748 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134248.10]
  assign _GEN_734 = _T_2838 ? 1'h0 : _GEN_504; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134249.10]
  assign _T_2839 = _T_2765 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134252.10]
  assign _GEN_735 = _T_2839 ? 1'h0 : _GEN_505; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134253.10]
  assign _GEN_736 = io_sfence_bits_rs2 & _GEN_732; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134099.8]
  assign _GEN_737 = io_sfence_bits_rs2 & _GEN_733; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134099.8]
  assign _GEN_738 = io_sfence_bits_rs2 & _GEN_734; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134099.8]
  assign _GEN_739 = io_sfence_bits_rs2 & _GEN_735; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134099.8]
  assign _T_2845 = _T_404[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@134272.8]
  assign _T_2846 = _T_2845 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@134273.8]
  assign _T_2849 = sectored_entries_4_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134280.10]
  assign _T_2861 = sectored_entries_4_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134304.10]
  assign _T_2866 = sectored_entries_4_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134315.10]
  assign _T_2878 = sectored_entries_4_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134339.10]
  assign _T_2883 = sectored_entries_4_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134350.10]
  assign _T_2895 = sectored_entries_4_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134374.10]
  assign _T_2900 = sectored_entries_4_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134385.10]
  assign _T_2912 = sectored_entries_4_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134409.10]
  assign _T_2983 = _T_2861 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134571.10]
  assign _GEN_760 = _T_2983 ? 1'h0 : _GEN_512; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134572.10]
  assign _T_2984 = _T_2878 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134575.10]
  assign _GEN_761 = _T_2984 ? 1'h0 : _GEN_513; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134576.10]
  assign _T_2985 = _T_2895 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134579.10]
  assign _GEN_762 = _T_2985 ? 1'h0 : _GEN_514; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134580.10]
  assign _T_2986 = _T_2912 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134583.10]
  assign _GEN_763 = _T_2986 ? 1'h0 : _GEN_515; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134584.10]
  assign _GEN_764 = io_sfence_bits_rs2 & _GEN_760; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134430.8]
  assign _GEN_765 = io_sfence_bits_rs2 & _GEN_761; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134430.8]
  assign _GEN_766 = io_sfence_bits_rs2 & _GEN_762; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134430.8]
  assign _GEN_767 = io_sfence_bits_rs2 & _GEN_763; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134430.8]
  assign _T_2992 = _T_410[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@134603.8]
  assign _T_2993 = _T_2992 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@134604.8]
  assign _T_2996 = sectored_entries_5_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134611.10]
  assign _T_3008 = sectored_entries_5_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134635.10]
  assign _T_3013 = sectored_entries_5_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134646.10]
  assign _T_3025 = sectored_entries_5_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134670.10]
  assign _T_3030 = sectored_entries_5_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134681.10]
  assign _T_3042 = sectored_entries_5_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134705.10]
  assign _T_3047 = sectored_entries_5_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134716.10]
  assign _T_3059 = sectored_entries_5_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134740.10]
  assign _T_3130 = _T_3008 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134902.10]
  assign _GEN_788 = _T_3130 ? 1'h0 : _GEN_522; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134903.10]
  assign _T_3131 = _T_3025 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134906.10]
  assign _GEN_789 = _T_3131 ? 1'h0 : _GEN_523; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134907.10]
  assign _T_3132 = _T_3042 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134910.10]
  assign _GEN_790 = _T_3132 ? 1'h0 : _GEN_524; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134911.10]
  assign _T_3133 = _T_3059 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@134914.10]
  assign _GEN_791 = _T_3133 ? 1'h0 : _GEN_525; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@134915.10]
  assign _GEN_792 = io_sfence_bits_rs2 & _GEN_788; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134761.8]
  assign _GEN_793 = io_sfence_bits_rs2 & _GEN_789; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134761.8]
  assign _GEN_794 = io_sfence_bits_rs2 & _GEN_790; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134761.8]
  assign _GEN_795 = io_sfence_bits_rs2 & _GEN_791; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@134761.8]
  assign _T_3139 = _T_416[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@134934.8]
  assign _T_3140 = _T_3139 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@134935.8]
  assign _T_3143 = sectored_entries_6_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134942.10]
  assign _T_3155 = sectored_entries_6_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134966.10]
  assign _T_3160 = sectored_entries_6_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@134977.10]
  assign _T_3172 = sectored_entries_6_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135001.10]
  assign _T_3177 = sectored_entries_6_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135012.10]
  assign _T_3189 = sectored_entries_6_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135036.10]
  assign _T_3194 = sectored_entries_6_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135047.10]
  assign _T_3206 = sectored_entries_6_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135071.10]
  assign _T_3277 = _T_3155 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135233.10]
  assign _GEN_816 = _T_3277 ? 1'h0 : _GEN_532; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135234.10]
  assign _T_3278 = _T_3172 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135237.10]
  assign _GEN_817 = _T_3278 ? 1'h0 : _GEN_533; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135238.10]
  assign _T_3279 = _T_3189 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135241.10]
  assign _GEN_818 = _T_3279 ? 1'h0 : _GEN_534; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135242.10]
  assign _T_3280 = _T_3206 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135245.10]
  assign _GEN_819 = _T_3280 ? 1'h0 : _GEN_535; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135246.10]
  assign _GEN_820 = io_sfence_bits_rs2 & _GEN_816; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135092.8]
  assign _GEN_821 = io_sfence_bits_rs2 & _GEN_817; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135092.8]
  assign _GEN_822 = io_sfence_bits_rs2 & _GEN_818; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135092.8]
  assign _GEN_823 = io_sfence_bits_rs2 & _GEN_819; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135092.8]
  assign _T_3286 = _T_422[19:10]; // @[TLB.scala 148:28:freechips.rocketchip.system.DefaultRV32Config.fir@135265.8]
  assign _T_3287 = _T_3286 == 10'h0; // @[TLB.scala 148:63:freechips.rocketchip.system.DefaultRV32Config.fir@135266.8]
  assign _T_3290 = sectored_entries_7_data_0[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135273.10]
  assign _T_3302 = sectored_entries_7_data_0[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135297.10]
  assign _T_3307 = sectored_entries_7_data_1[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135308.10]
  assign _T_3319 = sectored_entries_7_data_1[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135332.10]
  assign _T_3324 = sectored_entries_7_data_2[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135343.10]
  assign _T_3336 = sectored_entries_7_data_2[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135367.10]
  assign _T_3341 = sectored_entries_7_data_3[0]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135378.10]
  assign _T_3353 = sectored_entries_7_data_3[12]; // @[TLB.scala 96:41:freechips.rocketchip.system.DefaultRV32Config.fir@135402.10]
  assign _T_3424 = _T_3302 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135564.10]
  assign _GEN_844 = _T_3424 ? 1'h0 : _GEN_542; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135565.10]
  assign _T_3425 = _T_3319 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135568.10]
  assign _GEN_845 = _T_3425 ? 1'h0 : _GEN_543; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135569.10]
  assign _T_3426 = _T_3336 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135572.10]
  assign _GEN_846 = _T_3426 ? 1'h0 : _GEN_544; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135573.10]
  assign _T_3427 = _T_3353 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135576.10]
  assign _GEN_847 = _T_3427 ? 1'h0 : _GEN_545; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135577.10]
  assign _GEN_848 = io_sfence_bits_rs2 & _GEN_844; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135423.8]
  assign _GEN_849 = io_sfence_bits_rs2 & _GEN_845; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135423.8]
  assign _GEN_850 = io_sfence_bits_rs2 & _GEN_846; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135423.8]
  assign _GEN_851 = io_sfence_bits_rs2 & _GEN_847; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135423.8]
  assign _T_3459 = _T_758 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135643.10]
  assign _GEN_857 = _T_3459 ? 1'h0 : _GEN_458; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135644.10]
  assign _GEN_858 = io_sfence_bits_rs2 & _GEN_857; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135607.8]
  assign _T_3491 = _T_782 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135707.10]
  assign _GEN_861 = _T_3491 ? 1'h0 : _GEN_462; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135708.10]
  assign _GEN_862 = io_sfence_bits_rs2 & _GEN_861; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135671.8]
  assign _T_3523 = _T_806 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135771.10]
  assign _GEN_865 = _T_3523 ? 1'h0 : _GEN_466; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135772.10]
  assign _GEN_866 = io_sfence_bits_rs2 & _GEN_865; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135735.8]
  assign _T_3555 = _T_830 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135835.10]
  assign _GEN_869 = _T_3555 ? 1'h0 : _GEN_470; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135836.10]
  assign _GEN_870 = io_sfence_bits_rs2 & _GEN_869; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135799.8]
  assign _T_3587 = _T_21 == 1'h0; // @[TLB.scala 156:15:freechips.rocketchip.system.DefaultRV32Config.fir@135899.10]
  assign _GEN_873 = _T_3587 ? 1'h0 : _GEN_454; // @[TLB.scala 156:21:freechips.rocketchip.system.DefaultRV32Config.fir@135900.10]
  assign _GEN_874 = io_sfence_bits_rs2 & _GEN_873; // @[TLB.scala 371:40:freechips.rocketchip.system.DefaultRV32Config.fir@135863.8]
  assign _T_3589 = multipleHits | reset; // @[TLB.scala 375:24:freechips.rocketchip.system.DefaultRV32Config.fir@135909.4]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 324:16:freechips.rocketchip.system.DefaultRV32Config.fir@132717.4]
  assign io_resp_miss = _T_2107 | multipleHits; // @[TLB.scala 337:16:freechips.rocketchip.system.DefaultRV32Config.fir@132761.4]
  assign io_resp_paddr = {ppn,_T_33}; // @[TLB.scala 338:17:freechips.rocketchip.system.DefaultRV32Config.fir@132764.4]
  assign io_resp_pf_inst = _T_2086 != 14'h0; // @[TLB.scala 327:19:freechips.rocketchip.system.DefaultRV32Config.fir@132731.4]
  assign io_resp_ae_inst = _T_2094 != 14'h0; // @[TLB.scala 330:19:freechips.rocketchip.system.DefaultRV32Config.fir@132741.4]
  assign io_resp_cacheable = _T_2100 != 14'h0; // @[TLB.scala 334:21:freechips.rocketchip.system.DefaultRV32Config.fir@132751.4]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 340:20:freechips.rocketchip.system.DefaultRV32Config.fir@132766.4]
  assign io_ptw_req_bits_valid = io_kill == 1'h0; // @[TLB.scala 341:25:freechips.rocketchip.system.DefaultRV32Config.fir@132768.4]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 342:29:freechips.rocketchip.system.DefaultRV32Config.fir@132769.4]
  assign _2_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign _2_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@129524.4]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 193:14:freechips.rocketchip.system.DefaultRV32Config.fir@129555.4]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129547.4]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129547.4]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129547.4]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129547.4]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129547.4]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129547.4]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129547.4]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129548.4]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129548.4]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129548.4]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129548.4]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129548.4]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129548.4]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129548.4]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129549.4]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129549.4]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129549.4]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129549.4]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129549.4]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129549.4]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129549.4]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129550.4]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129550.4]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129550.4]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129550.4]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129550.4]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129550.4]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129550.4]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129551.4]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129551.4]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129551.4]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129551.4]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129551.4]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129551.4]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129551.4]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129552.4]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129552.4]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129552.4]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129552.4]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129552.4]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129552.4]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129552.4]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129553.4]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129553.4]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129553.4]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129553.4]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129553.4]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129553.4]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129553.4]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129554.4]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129554.4]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129554.4]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129554.4]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129554.4]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129554.4]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 192:14:freechips.rocketchip.system.DefaultRV32Config.fir@129554.4]
  assign pmp_io_addr = {mpu_ppn,_T_33}; // @[TLB.scala 190:15:freechips.rocketchip.system.DefaultRV32Config.fir@129545.4]
  assign _2_1_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_u = _GEN_35[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_px = _GEN_35[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_1_io_x_c = _GEN_35[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130210.4]
  assign _2_2_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_u = _GEN_39[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_px = _GEN_39[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_2_io_x_c = _GEN_39[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130251.4]
  assign _2_3_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_u = _GEN_43[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_px = _GEN_43[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_3_io_x_c = _GEN_43[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130292.4]
  assign _2_4_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_u = _GEN_47[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_px = _GEN_47[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_4_io_x_c = _GEN_47[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130333.4]
  assign _2_5_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_u = _GEN_51[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_px = _GEN_51[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_5_io_x_c = _GEN_51[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130374.4]
  assign _2_6_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_u = _GEN_55[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_px = _GEN_55[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_6_io_x_c = _GEN_55[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130415.4]
  assign _2_7_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_u = _GEN_59[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_px = _GEN_59[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_7_io_x_c = _GEN_59[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130456.4]
  assign _2_8_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_u = _GEN_63[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_px = _GEN_63[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_8_io_x_c = _GEN_63[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130497.4]
  assign _2_9_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_9_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130537.4]
  assign _2_10_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_10_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130584.4]
  assign _2_11_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_11_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130631.4]
  assign _2_12_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_12_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130678.4]
  assign _2_13_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_13_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@130725.4]
  assign _2_14_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_u = _GEN_35[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_px = _GEN_35[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_14_io_x_c = _GEN_35[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131190.4]
  assign _2_15_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_u = _GEN_39[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_px = _GEN_39[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_15_io_x_c = _GEN_39[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131231.4]
  assign _2_16_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_u = _GEN_43[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_px = _GEN_43[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_16_io_x_c = _GEN_43[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131272.4]
  assign _2_17_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_u = _GEN_47[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_px = _GEN_47[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_17_io_x_c = _GEN_47[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131313.4]
  assign _2_18_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_u = _GEN_51[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_px = _GEN_51[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_18_io_x_c = _GEN_51[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131354.4]
  assign _2_19_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_u = _GEN_55[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_px = _GEN_55[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_19_io_x_c = _GEN_55[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131395.4]
  assign _2_20_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_u = _GEN_59[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_px = _GEN_59[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_20_io_x_c = _GEN_59[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131436.4]
  assign _2_21_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_u = _GEN_63[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_px = _GEN_63[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_21_io_x_c = _GEN_63[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131477.4]
  assign _2_22_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_22_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131517.4]
  assign _2_23_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_23_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131557.4]
  assign _2_24_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_24_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131597.4]
  assign _2_25_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_25_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131637.4]
  assign _2_26_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_26_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131677.4]
  assign _2_27_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_u = _GEN_35[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_px = _GEN_35[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_27_io_x_c = _GEN_35[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131718.4]
  assign _2_28_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_u = _GEN_39[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_px = _GEN_39[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_28_io_x_c = _GEN_39[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131759.4]
  assign _2_29_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_u = _GEN_43[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_px = _GEN_43[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_29_io_x_c = _GEN_43[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131800.4]
  assign _2_30_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_u = _GEN_47[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_px = _GEN_47[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_30_io_x_c = _GEN_47[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131841.4]
  assign _2_31_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_u = _GEN_51[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_px = _GEN_51[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_31_io_x_c = _GEN_51[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131882.4]
  assign _2_32_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_u = _GEN_55[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_px = _GEN_55[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_32_io_x_c = _GEN_55[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131923.4]
  assign _2_33_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_u = _GEN_59[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_px = _GEN_59[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_33_io_x_c = _GEN_59[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@131964.4]
  assign _2_34_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_u = _GEN_63[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_px = _GEN_63[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_34_io_x_c = _GEN_63[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132005.4]
  assign _2_35_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_35_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132045.4]
  assign _2_36_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_36_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132085.4]
  assign _2_37_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_37_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132125.4]
  assign _2_38_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
  assign _2_38_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:freechips.rocketchip.system.DefaultRV32Config.fir@132165.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_72[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_73[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_75[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_76[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_78[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_79[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_81[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_82[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  special_entry_level = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  special_entry_tag = _RAND_85[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_86[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  state = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  r_refill_tag = _RAND_89[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_90[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_92[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_sectored_hit = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1904 = _RAND_94[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1905 = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            sectored_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            if (2'h0 == _T_996) begin
              sectored_entries_0_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            if (2'h1 == _T_996) begin
              sectored_entries_0_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            if (2'h2 == _T_996) begin
              sectored_entries_0_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_994) begin
            if (2'h3 == _T_996) begin
              sectored_entries_0_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2258) begin
            if (_T_2261) begin
              sectored_entries_0_valid_0 <= 1'h0;
            end else begin
              if (_T_382) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_0_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_994) begin
                          sectored_entries_0_valid_0 <= _GEN_84;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_0 <= _GEN_84;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_382) begin
              if (2'h0 == _T_477) begin
                sectored_entries_0_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_0 <= _GEN_84;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_994) begin
                      sectored_entries_0_valid_0 <= _GEN_84;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_0_valid_0 <= _GEN_652;
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_472;
      end
    end
    if (_T_3589) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2258) begin
            if (_T_2278) begin
              sectored_entries_0_valid_1 <= 1'h0;
            end else begin
              if (_T_382) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_0_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_994) begin
                          sectored_entries_0_valid_1 <= _GEN_85;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_1 <= _GEN_85;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_382) begin
              if (2'h1 == _T_477) begin
                sectored_entries_0_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_1 <= _GEN_85;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_994) begin
                      sectored_entries_0_valid_1 <= _GEN_85;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_0_valid_1 <= _GEN_653;
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_473;
      end
    end
    if (_T_3589) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2258) begin
            if (_T_2295) begin
              sectored_entries_0_valid_2 <= 1'h0;
            end else begin
              if (_T_382) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_0_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_994) begin
                          sectored_entries_0_valid_2 <= _GEN_86;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_2 <= _GEN_86;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_382) begin
              if (2'h2 == _T_477) begin
                sectored_entries_0_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_2 <= _GEN_86;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_994) begin
                      sectored_entries_0_valid_2 <= _GEN_86;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_0_valid_2 <= _GEN_654;
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_474;
      end
    end
    if (_T_3589) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2258) begin
            if (_T_2312) begin
              sectored_entries_0_valid_3 <= 1'h0;
            end else begin
              if (_T_382) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_0_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_994) begin
                          sectored_entries_0_valid_3 <= _GEN_87;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_3 <= _GEN_87;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_382) begin
              if (2'h3 == _T_477) begin
                sectored_entries_0_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_994) begin
                        sectored_entries_0_valid_3 <= _GEN_87;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_994) begin
                      sectored_entries_0_valid_3 <= _GEN_87;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_0_valid_3 <= _GEN_655;
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_475;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            sectored_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            if (2'h0 == _T_996) begin
              sectored_entries_1_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            if (2'h1 == _T_996) begin
              sectored_entries_1_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            if (2'h2 == _T_996) begin
              sectored_entries_1_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1011) begin
            if (2'h3 == _T_996) begin
              sectored_entries_1_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2405) begin
            if (_T_2408) begin
              sectored_entries_1_valid_0 <= 1'h0;
            end else begin
              if (_T_388) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_1_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1011) begin
                          sectored_entries_1_valid_0 <= _GEN_106;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_0 <= _GEN_106;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_388) begin
              if (2'h0 == _T_477) begin
                sectored_entries_1_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_0 <= _GEN_106;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1011) begin
                      sectored_entries_1_valid_0 <= _GEN_106;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_1_valid_0 <= _GEN_680;
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_482;
      end
    end
    if (_T_3589) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2405) begin
            if (_T_2425) begin
              sectored_entries_1_valid_1 <= 1'h0;
            end else begin
              if (_T_388) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_1_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1011) begin
                          sectored_entries_1_valid_1 <= _GEN_107;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_1 <= _GEN_107;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_388) begin
              if (2'h1 == _T_477) begin
                sectored_entries_1_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_1 <= _GEN_107;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1011) begin
                      sectored_entries_1_valid_1 <= _GEN_107;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_1_valid_1 <= _GEN_681;
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_483;
      end
    end
    if (_T_3589) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2405) begin
            if (_T_2442) begin
              sectored_entries_1_valid_2 <= 1'h0;
            end else begin
              if (_T_388) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_1_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1011) begin
                          sectored_entries_1_valid_2 <= _GEN_108;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_2 <= _GEN_108;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_388) begin
              if (2'h2 == _T_477) begin
                sectored_entries_1_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_2 <= _GEN_108;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1011) begin
                      sectored_entries_1_valid_2 <= _GEN_108;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_1_valid_2 <= _GEN_682;
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_484;
      end
    end
    if (_T_3589) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2405) begin
            if (_T_2459) begin
              sectored_entries_1_valid_3 <= 1'h0;
            end else begin
              if (_T_388) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_1_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1011) begin
                          sectored_entries_1_valid_3 <= _GEN_109;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_3 <= _GEN_109;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_388) begin
              if (2'h3 == _T_477) begin
                sectored_entries_1_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1011) begin
                        sectored_entries_1_valid_3 <= _GEN_109;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1011) begin
                      sectored_entries_1_valid_3 <= _GEN_109;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_1_valid_3 <= _GEN_683;
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_485;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            sectored_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            if (2'h0 == _T_996) begin
              sectored_entries_2_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            if (2'h1 == _T_996) begin
              sectored_entries_2_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            if (2'h2 == _T_996) begin
              sectored_entries_2_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1028) begin
            if (2'h3 == _T_996) begin
              sectored_entries_2_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2552) begin
            if (_T_2555) begin
              sectored_entries_2_valid_0 <= 1'h0;
            end else begin
              if (_T_394) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_2_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1028) begin
                          sectored_entries_2_valid_0 <= _GEN_128;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_0 <= _GEN_128;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_394) begin
              if (2'h0 == _T_477) begin
                sectored_entries_2_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_0 <= _GEN_128;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1028) begin
                      sectored_entries_2_valid_0 <= _GEN_128;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_2_valid_0 <= _GEN_708;
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_492;
      end
    end
    if (_T_3589) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2552) begin
            if (_T_2572) begin
              sectored_entries_2_valid_1 <= 1'h0;
            end else begin
              if (_T_394) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_2_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1028) begin
                          sectored_entries_2_valid_1 <= _GEN_129;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_1 <= _GEN_129;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_394) begin
              if (2'h1 == _T_477) begin
                sectored_entries_2_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_1 <= _GEN_129;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1028) begin
                      sectored_entries_2_valid_1 <= _GEN_129;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_2_valid_1 <= _GEN_709;
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_493;
      end
    end
    if (_T_3589) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2552) begin
            if (_T_2589) begin
              sectored_entries_2_valid_2 <= 1'h0;
            end else begin
              if (_T_394) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_2_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1028) begin
                          sectored_entries_2_valid_2 <= _GEN_130;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_2 <= _GEN_130;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_394) begin
              if (2'h2 == _T_477) begin
                sectored_entries_2_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_2 <= _GEN_130;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1028) begin
                      sectored_entries_2_valid_2 <= _GEN_130;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_2_valid_2 <= _GEN_710;
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_494;
      end
    end
    if (_T_3589) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2552) begin
            if (_T_2606) begin
              sectored_entries_2_valid_3 <= 1'h0;
            end else begin
              if (_T_394) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_2_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1028) begin
                          sectored_entries_2_valid_3 <= _GEN_131;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_3 <= _GEN_131;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_394) begin
              if (2'h3 == _T_477) begin
                sectored_entries_2_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1028) begin
                        sectored_entries_2_valid_3 <= _GEN_131;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1028) begin
                      sectored_entries_2_valid_3 <= _GEN_131;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_2_valid_3 <= _GEN_711;
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_495;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            sectored_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            if (2'h0 == _T_996) begin
              sectored_entries_3_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            if (2'h1 == _T_996) begin
              sectored_entries_3_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            if (2'h2 == _T_996) begin
              sectored_entries_3_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1045) begin
            if (2'h3 == _T_996) begin
              sectored_entries_3_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2699) begin
            if (_T_2702) begin
              sectored_entries_3_valid_0 <= 1'h0;
            end else begin
              if (_T_400) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_3_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1045) begin
                          sectored_entries_3_valid_0 <= _GEN_150;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_0 <= _GEN_150;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_400) begin
              if (2'h0 == _T_477) begin
                sectored_entries_3_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_0 <= _GEN_150;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1045) begin
                      sectored_entries_3_valid_0 <= _GEN_150;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_3_valid_0 <= _GEN_736;
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_502;
      end
    end
    if (_T_3589) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2699) begin
            if (_T_2719) begin
              sectored_entries_3_valid_1 <= 1'h0;
            end else begin
              if (_T_400) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_3_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1045) begin
                          sectored_entries_3_valid_1 <= _GEN_151;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_1 <= _GEN_151;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_400) begin
              if (2'h1 == _T_477) begin
                sectored_entries_3_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_1 <= _GEN_151;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1045) begin
                      sectored_entries_3_valid_1 <= _GEN_151;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_3_valid_1 <= _GEN_737;
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_503;
      end
    end
    if (_T_3589) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2699) begin
            if (_T_2736) begin
              sectored_entries_3_valid_2 <= 1'h0;
            end else begin
              if (_T_400) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_3_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1045) begin
                          sectored_entries_3_valid_2 <= _GEN_152;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_2 <= _GEN_152;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_400) begin
              if (2'h2 == _T_477) begin
                sectored_entries_3_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_2 <= _GEN_152;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1045) begin
                      sectored_entries_3_valid_2 <= _GEN_152;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_3_valid_2 <= _GEN_738;
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_504;
      end
    end
    if (_T_3589) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2699) begin
            if (_T_2753) begin
              sectored_entries_3_valid_3 <= 1'h0;
            end else begin
              if (_T_400) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_3_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1045) begin
                          sectored_entries_3_valid_3 <= _GEN_153;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_3 <= _GEN_153;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_400) begin
              if (2'h3 == _T_477) begin
                sectored_entries_3_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1045) begin
                        sectored_entries_3_valid_3 <= _GEN_153;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1045) begin
                      sectored_entries_3_valid_3 <= _GEN_153;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_3_valid_3 <= _GEN_739;
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_505;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            sectored_entries_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            if (2'h0 == _T_996) begin
              sectored_entries_4_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            if (2'h1 == _T_996) begin
              sectored_entries_4_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            if (2'h2 == _T_996) begin
              sectored_entries_4_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1062) begin
            if (2'h3 == _T_996) begin
              sectored_entries_4_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2846) begin
            if (_T_2849) begin
              sectored_entries_4_valid_0 <= 1'h0;
            end else begin
              if (_T_406) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_4_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1062) begin
                          sectored_entries_4_valid_0 <= _GEN_172;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_0 <= _GEN_172;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_406) begin
              if (2'h0 == _T_477) begin
                sectored_entries_4_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_0 <= _GEN_172;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1062) begin
                      sectored_entries_4_valid_0 <= _GEN_172;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_4_valid_0 <= _GEN_764;
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_512;
      end
    end
    if (_T_3589) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2846) begin
            if (_T_2866) begin
              sectored_entries_4_valid_1 <= 1'h0;
            end else begin
              if (_T_406) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_4_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1062) begin
                          sectored_entries_4_valid_1 <= _GEN_173;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_1 <= _GEN_173;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_406) begin
              if (2'h1 == _T_477) begin
                sectored_entries_4_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_1 <= _GEN_173;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1062) begin
                      sectored_entries_4_valid_1 <= _GEN_173;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_4_valid_1 <= _GEN_765;
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_513;
      end
    end
    if (_T_3589) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2846) begin
            if (_T_2883) begin
              sectored_entries_4_valid_2 <= 1'h0;
            end else begin
              if (_T_406) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_4_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1062) begin
                          sectored_entries_4_valid_2 <= _GEN_174;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_2 <= _GEN_174;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_406) begin
              if (2'h2 == _T_477) begin
                sectored_entries_4_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_2 <= _GEN_174;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1062) begin
                      sectored_entries_4_valid_2 <= _GEN_174;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_4_valid_2 <= _GEN_766;
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_514;
      end
    end
    if (_T_3589) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2846) begin
            if (_T_2900) begin
              sectored_entries_4_valid_3 <= 1'h0;
            end else begin
              if (_T_406) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_4_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1062) begin
                          sectored_entries_4_valid_3 <= _GEN_175;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_3 <= _GEN_175;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_406) begin
              if (2'h3 == _T_477) begin
                sectored_entries_4_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1062) begin
                        sectored_entries_4_valid_3 <= _GEN_175;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1062) begin
                      sectored_entries_4_valid_3 <= _GEN_175;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_4_valid_3 <= _GEN_767;
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_515;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            sectored_entries_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            if (2'h0 == _T_996) begin
              sectored_entries_5_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            if (2'h1 == _T_996) begin
              sectored_entries_5_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            if (2'h2 == _T_996) begin
              sectored_entries_5_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1079) begin
            if (2'h3 == _T_996) begin
              sectored_entries_5_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2993) begin
            if (_T_2996) begin
              sectored_entries_5_valid_0 <= 1'h0;
            end else begin
              if (_T_412) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_5_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1079) begin
                          sectored_entries_5_valid_0 <= _GEN_194;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_0 <= _GEN_194;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_412) begin
              if (2'h0 == _T_477) begin
                sectored_entries_5_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_0 <= _GEN_194;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1079) begin
                      sectored_entries_5_valid_0 <= _GEN_194;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_5_valid_0 <= _GEN_792;
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_522;
      end
    end
    if (_T_3589) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2993) begin
            if (_T_3013) begin
              sectored_entries_5_valid_1 <= 1'h0;
            end else begin
              if (_T_412) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_5_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1079) begin
                          sectored_entries_5_valid_1 <= _GEN_195;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_1 <= _GEN_195;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_412) begin
              if (2'h1 == _T_477) begin
                sectored_entries_5_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_1 <= _GEN_195;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1079) begin
                      sectored_entries_5_valid_1 <= _GEN_195;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_5_valid_1 <= _GEN_793;
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_523;
      end
    end
    if (_T_3589) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2993) begin
            if (_T_3030) begin
              sectored_entries_5_valid_2 <= 1'h0;
            end else begin
              if (_T_412) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_5_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1079) begin
                          sectored_entries_5_valid_2 <= _GEN_196;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_2 <= _GEN_196;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_412) begin
              if (2'h2 == _T_477) begin
                sectored_entries_5_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_2 <= _GEN_196;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1079) begin
                      sectored_entries_5_valid_2 <= _GEN_196;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_5_valid_2 <= _GEN_794;
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_524;
      end
    end
    if (_T_3589) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_2993) begin
            if (_T_3047) begin
              sectored_entries_5_valid_3 <= 1'h0;
            end else begin
              if (_T_412) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_5_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1079) begin
                          sectored_entries_5_valid_3 <= _GEN_197;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_3 <= _GEN_197;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_412) begin
              if (2'h3 == _T_477) begin
                sectored_entries_5_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1079) begin
                        sectored_entries_5_valid_3 <= _GEN_197;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1079) begin
                      sectored_entries_5_valid_3 <= _GEN_197;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_5_valid_3 <= _GEN_795;
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_525;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            sectored_entries_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            if (2'h0 == _T_996) begin
              sectored_entries_6_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            if (2'h1 == _T_996) begin
              sectored_entries_6_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            if (2'h2 == _T_996) begin
              sectored_entries_6_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1096) begin
            if (2'h3 == _T_996) begin
              sectored_entries_6_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3140) begin
            if (_T_3143) begin
              sectored_entries_6_valid_0 <= 1'h0;
            end else begin
              if (_T_418) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_6_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1096) begin
                          sectored_entries_6_valid_0 <= _GEN_216;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_0 <= _GEN_216;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_418) begin
              if (2'h0 == _T_477) begin
                sectored_entries_6_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_0 <= _GEN_216;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1096) begin
                      sectored_entries_6_valid_0 <= _GEN_216;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_6_valid_0 <= _GEN_820;
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_532;
      end
    end
    if (_T_3589) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3140) begin
            if (_T_3160) begin
              sectored_entries_6_valid_1 <= 1'h0;
            end else begin
              if (_T_418) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_6_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1096) begin
                          sectored_entries_6_valid_1 <= _GEN_217;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_1 <= _GEN_217;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_418) begin
              if (2'h1 == _T_477) begin
                sectored_entries_6_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_1 <= _GEN_217;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1096) begin
                      sectored_entries_6_valid_1 <= _GEN_217;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_6_valid_1 <= _GEN_821;
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_533;
      end
    end
    if (_T_3589) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3140) begin
            if (_T_3177) begin
              sectored_entries_6_valid_2 <= 1'h0;
            end else begin
              if (_T_418) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_6_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1096) begin
                          sectored_entries_6_valid_2 <= _GEN_218;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_2 <= _GEN_218;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_418) begin
              if (2'h2 == _T_477) begin
                sectored_entries_6_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_2 <= _GEN_218;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1096) begin
                      sectored_entries_6_valid_2 <= _GEN_218;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_6_valid_2 <= _GEN_822;
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_534;
      end
    end
    if (_T_3589) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3140) begin
            if (_T_3194) begin
              sectored_entries_6_valid_3 <= 1'h0;
            end else begin
              if (_T_418) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_6_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1096) begin
                          sectored_entries_6_valid_3 <= _GEN_219;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_3 <= _GEN_219;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_418) begin
              if (2'h3 == _T_477) begin
                sectored_entries_6_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1096) begin
                        sectored_entries_6_valid_3 <= _GEN_219;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1096) begin
                      sectored_entries_6_valid_3 <= _GEN_219;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_6_valid_3 <= _GEN_823;
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_535;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            sectored_entries_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            if (2'h0 == _T_996) begin
              sectored_entries_7_data_0 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            if (2'h1 == _T_996) begin
              sectored_entries_7_data_1 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            if (2'h2 == _T_996) begin
              sectored_entries_7_data_2 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (!(_T_932)) begin
          if (_T_1113) begin
            if (2'h3 == _T_996) begin
              sectored_entries_7_data_3 <= _T_931;
            end
          end
        end
      end
    end
    if (_T_3589) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3287) begin
            if (_T_3290) begin
              sectored_entries_7_valid_0 <= 1'h0;
            end else begin
              if (_T_424) begin
                if (2'h0 == _T_477) begin
                  sectored_entries_7_valid_0 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1113) begin
                          sectored_entries_7_valid_0 <= _GEN_238;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_0 <= _GEN_238;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_424) begin
              if (2'h0 == _T_477) begin
                sectored_entries_7_valid_0 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_0 <= _GEN_238;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1113) begin
                      sectored_entries_7_valid_0 <= _GEN_238;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_7_valid_0 <= _GEN_848;
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_542;
      end
    end
    if (_T_3589) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3287) begin
            if (_T_3307) begin
              sectored_entries_7_valid_1 <= 1'h0;
            end else begin
              if (_T_424) begin
                if (2'h1 == _T_477) begin
                  sectored_entries_7_valid_1 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1113) begin
                          sectored_entries_7_valid_1 <= _GEN_239;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_1 <= _GEN_239;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_424) begin
              if (2'h1 == _T_477) begin
                sectored_entries_7_valid_1 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_1 <= _GEN_239;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1113) begin
                      sectored_entries_7_valid_1 <= _GEN_239;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_7_valid_1 <= _GEN_849;
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_543;
      end
    end
    if (_T_3589) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3287) begin
            if (_T_3324) begin
              sectored_entries_7_valid_2 <= 1'h0;
            end else begin
              if (_T_424) begin
                if (2'h2 == _T_477) begin
                  sectored_entries_7_valid_2 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1113) begin
                          sectored_entries_7_valid_2 <= _GEN_240;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_2 <= _GEN_240;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_424) begin
              if (2'h2 == _T_477) begin
                sectored_entries_7_valid_2 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_2 <= _GEN_240;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1113) begin
                      sectored_entries_7_valid_2 <= _GEN_240;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_7_valid_2 <= _GEN_850;
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_544;
      end
    end
    if (_T_3589) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_3287) begin
            if (_T_3341) begin
              sectored_entries_7_valid_3 <= 1'h0;
            end else begin
              if (_T_424) begin
                if (2'h3 == _T_477) begin
                  sectored_entries_7_valid_3 <= 1'h0;
                end else begin
                  if (_T_893) begin
                    if (!(_T_915)) begin
                      if (!(_T_932)) begin
                        if (_T_1113) begin
                          sectored_entries_7_valid_3 <= _GEN_241;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_3 <= _GEN_241;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_424) begin
              if (2'h3 == _T_477) begin
                sectored_entries_7_valid_3 <= 1'h0;
              end else begin
                if (_T_893) begin
                  if (!(_T_915)) begin
                    if (!(_T_932)) begin
                      if (_T_1113) begin
                        sectored_entries_7_valid_3 <= _GEN_241;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_893) begin
                if (!(_T_915)) begin
                  if (!(_T_932)) begin
                    if (_T_1113) begin
                      sectored_entries_7_valid_3 <= _GEN_241;
                    end
                  end
                end
              end
            end
          end
        end else begin
          sectored_entries_7_valid_3 <= _GEN_851;
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_545;
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_933) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_933) begin
            superpage_entries_0_data_0 <= _T_931;
          end
        end
      end
    end
    if (_T_3589) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (superpage_hits_0) begin
            superpage_entries_0_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              if (!(_T_915)) begin
                if (_T_932) begin
                  superpage_entries_0_valid_0 <= _GEN_66;
                end
              end
            end
          end
        end else begin
          superpage_entries_0_valid_0 <= _GEN_858;
        end
      end else begin
        if (_T_893) begin
          if (!(_T_915)) begin
            if (_T_932) begin
              superpage_entries_0_valid_0 <= _GEN_66;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_948) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_948) begin
            superpage_entries_1_data_0 <= _T_931;
          end
        end
      end
    end
    if (_T_3589) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (superpage_hits_1) begin
            superpage_entries_1_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              if (!(_T_915)) begin
                if (_T_932) begin
                  superpage_entries_1_valid_0 <= _GEN_70;
                end
              end
            end
          end
        end else begin
          superpage_entries_1_valid_0 <= _GEN_862;
        end
      end else begin
        if (_T_893) begin
          if (!(_T_915)) begin
            if (_T_932) begin
              superpage_entries_1_valid_0 <= _GEN_70;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_963) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_963) begin
            superpage_entries_2_data_0 <= _T_931;
          end
        end
      end
    end
    if (_T_3589) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (superpage_hits_2) begin
            superpage_entries_2_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              if (!(_T_915)) begin
                if (_T_932) begin
                  superpage_entries_2_valid_0 <= _GEN_74;
                end
              end
            end
          end
        end else begin
          superpage_entries_2_valid_0 <= _GEN_866;
        end
      end else begin
        if (_T_893) begin
          if (!(_T_915)) begin
            if (_T_932) begin
              superpage_entries_2_valid_0 <= _GEN_74;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_978) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_893) begin
      if (!(_T_915)) begin
        if (_T_932) begin
          if (_T_978) begin
            superpage_entries_3_data_0 <= _T_931;
          end
        end
      end
    end
    if (_T_3589) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (superpage_hits_3) begin
            superpage_entries_3_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              if (!(_T_915)) begin
                if (_T_932) begin
                  superpage_entries_3_valid_0 <= _GEN_78;
                end
              end
            end
          end
        end else begin
          superpage_entries_3_valid_0 <= _GEN_870;
        end
      end else begin
        if (_T_893) begin
          if (!(_T_915)) begin
            if (_T_932) begin
              superpage_entries_3_valid_0 <= _GEN_78;
            end
          end
        end
      end
    end
    if (_T_893) begin
      if (_T_915) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (_T_893) begin
      if (_T_915) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (_T_893) begin
      if (_T_915) begin
        special_entry_data_0 <= _T_931;
      end
    end
    if (_T_3589) begin
      special_entry_valid_0 <= 1'h0;
    end else begin
      if (io_sfence_valid) begin
        if (io_sfence_bits_rs1) begin
          if (_T_586) begin
            special_entry_valid_0 <= 1'h0;
          end else begin
            if (_T_893) begin
              special_entry_valid_0 <= _GEN_354;
            end
          end
        end else begin
          special_entry_valid_0 <= _GEN_874;
        end
      end else begin
        if (_T_893) begin
          special_entry_valid_0 <= _GEN_354;
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (io_ptw_resp_valid) begin
        state <= 2'h0;
      end else begin
        if (_T_2244) begin
          state <= 2'h3;
        end else begin
          if (_T_4) begin
            if (io_kill) begin
              state <= 2'h0;
            end else begin
              if (io_ptw_req_ready) begin
                if (io_sfence_valid) begin
                  state <= 2'h3;
                end else begin
                  state <= 2'h2;
                end
              end else begin
                if (io_sfence_valid) begin
                  state <= 2'h0;
                end else begin
                  if (_T_2114) begin
                    state <= 2'h1;
                  end
                end
              end
            end
          end else begin
            if (_T_2114) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if (_T_2114) begin
      r_refill_tag <= vpn;
    end
    if (_T_2114) begin
      if (_T_2134) begin
        r_superpage_repl_addr <= _T_2130;
      end else begin
        if (_T_2136) begin
          r_superpage_repl_addr <= 2'h0;
        end else begin
          if (_T_2137) begin
            r_superpage_repl_addr <= 2'h1;
          end else begin
            if (_T_2138) begin
              r_superpage_repl_addr <= 2'h2;
            end else begin
              r_superpage_repl_addr <= 2'h3;
            end
          end
        end
      end
    end
    if (_T_2114) begin
      if (_T_2198) begin
        r_sectored_repl_addr <= _T_2166;
      end else begin
        if (_T_2200) begin
          r_sectored_repl_addr <= 3'h0;
        end else begin
          if (_T_2201) begin
            r_sectored_repl_addr <= 3'h1;
          end else begin
            if (_T_2202) begin
              r_sectored_repl_addr <= 3'h2;
            end else begin
              if (_T_2203) begin
                r_sectored_repl_addr <= 3'h3;
              end else begin
                if (_T_2204) begin
                  r_sectored_repl_addr <= 3'h4;
                end else begin
                  if (_T_2205) begin
                    r_sectored_repl_addr <= 3'h5;
                  end else begin
                    if (_T_2206) begin
                      r_sectored_repl_addr <= 3'h6;
                    end else begin
                      r_sectored_repl_addr <= 3'h7;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_2114) begin
      r_sectored_hit_addr <= _T_1931;
    end
    if (_T_2114) begin
      r_sectored_hit <= _T_1913;
    end
    if (_T_1906) begin
      if (_T_1913) begin
        _T_1904 <= _T_1960;
      end
    end
    if (_T_1906) begin
      if (_T_1963) begin
        _T_1905 <= _T_1992;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & _T_2251) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:368 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@132936.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & _T_2251) begin
          $fatal; // @[TLB.scala 368:13:freechips.rocketchip.system.DefaultRV32Config.fir@132937.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
`endif __TLB_1

