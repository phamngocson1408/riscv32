module RoundAnyRawFNToRecFN( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190939.2]
  input         io_invalidExc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  input         io_infiniteExc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  input         io_in_isNaN, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  input         io_in_isInf, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  input         io_in_isZero, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  input         io_in_sign, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  input  [9:0]  io_in_sExp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  input  [26:0] io_in_sig, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  input  [2:0]  io_roundingMode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  output [32:0] io_out, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
  output [4:0]  io_exceptionFlags // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190940.4]
);
  wire [8:0] my_lowMask_io_in; // @[RoundAnyRawFNToRecFN.scala 160:40:freechips.rocketchip.system.DefaultRV32Config.fir@190967.4]
  wire [24:0] my_lowMask_io_out; // @[RoundAnyRawFNToRecFN.scala 160:40:freechips.rocketchip.system.DefaultRV32Config.fir@190967.4]
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53:freechips.rocketchip.system.DefaultRV32Config.fir@190943.4]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53:freechips.rocketchip.system.DefaultRV32Config.fir@190945.4]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53:freechips.rocketchip.system.DefaultRV32Config.fir@190946.4]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53:freechips.rocketchip.system.DefaultRV32Config.fir@190947.4]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53:freechips.rocketchip.system.DefaultRV32Config.fir@190948.4]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27:freechips.rocketchip.system.DefaultRV32Config.fir@190949.4]
  wire  _T_1; // @[RoundAnyRawFNToRecFN.scala 96:66:freechips.rocketchip.system.DefaultRV32Config.fir@190950.4]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63:freechips.rocketchip.system.DefaultRV32Config.fir@190951.4]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42:freechips.rocketchip.system.DefaultRV32Config.fir@190952.4]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 120:61:freechips.rocketchip.system.DefaultRV32Config.fir@190954.4]
  wire [24:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 163:21:freechips.rocketchip.system.DefaultRV32Config.fir@190971.4]
  wire [24:0] _T_4; // @[RoundAnyRawFNToRecFN.scala 163:21:freechips.rocketchip.system.DefaultRV32Config.fir@190971.4]
  wire [26:0] roundMask; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190972.4]
  wire [26:0] shiftedRoundMask; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190974.4]
  wire [26:0] _T_6; // @[RoundAnyRawFNToRecFN.scala 170:28:freechips.rocketchip.system.DefaultRV32Config.fir@190975.4]
  wire [26:0] roundPosMask; // @[RoundAnyRawFNToRecFN.scala 170:46:freechips.rocketchip.system.DefaultRV32Config.fir@190976.4]
  wire [26:0] _T_7; // @[RoundAnyRawFNToRecFN.scala 172:40:freechips.rocketchip.system.DefaultRV32Config.fir@190977.4]
  wire  roundPosBit; // @[RoundAnyRawFNToRecFN.scala 172:56:freechips.rocketchip.system.DefaultRV32Config.fir@190978.4]
  wire [26:0] _T_8; // @[RoundAnyRawFNToRecFN.scala 174:42:freechips.rocketchip.system.DefaultRV32Config.fir@190979.4]
  wire  anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 174:62:freechips.rocketchip.system.DefaultRV32Config.fir@190980.4]
  wire  anyRound; // @[RoundAnyRawFNToRecFN.scala 176:36:freechips.rocketchip.system.DefaultRV32Config.fir@190981.4]
  wire  _T_9; // @[RoundAnyRawFNToRecFN.scala 180:38:freechips.rocketchip.system.DefaultRV32Config.fir@190982.4]
  wire  _T_10; // @[RoundAnyRawFNToRecFN.scala 180:67:freechips.rocketchip.system.DefaultRV32Config.fir@190983.4]
  wire  _T_11; // @[RoundAnyRawFNToRecFN.scala 182:29:freechips.rocketchip.system.DefaultRV32Config.fir@190984.4]
  wire  roundIncr; // @[RoundAnyRawFNToRecFN.scala 181:31:freechips.rocketchip.system.DefaultRV32Config.fir@190985.4]
  wire [26:0] _T_12; // @[RoundAnyRawFNToRecFN.scala 186:32:freechips.rocketchip.system.DefaultRV32Config.fir@190986.4]
  wire [25:0] _T_14; // @[RoundAnyRawFNToRecFN.scala 186:49:freechips.rocketchip.system.DefaultRV32Config.fir@190988.4]
  wire  _T_15; // @[RoundAnyRawFNToRecFN.scala 187:49:freechips.rocketchip.system.DefaultRV32Config.fir@190989.4]
  wire  _T_16; // @[RoundAnyRawFNToRecFN.scala 188:30:freechips.rocketchip.system.DefaultRV32Config.fir@190990.4]
  wire  _T_17; // @[RoundAnyRawFNToRecFN.scala 187:64:freechips.rocketchip.system.DefaultRV32Config.fir@190991.4]
  wire [25:0] _T_19; // @[RoundAnyRawFNToRecFN.scala 187:25:freechips.rocketchip.system.DefaultRV32Config.fir@190993.4]
  wire [25:0] _T_20; // @[RoundAnyRawFNToRecFN.scala 187:21:freechips.rocketchip.system.DefaultRV32Config.fir@190994.4]
  wire [25:0] _T_21; // @[RoundAnyRawFNToRecFN.scala 186:61:freechips.rocketchip.system.DefaultRV32Config.fir@190995.4]
  wire [26:0] _T_22; // @[RoundAnyRawFNToRecFN.scala 192:32:freechips.rocketchip.system.DefaultRV32Config.fir@190996.4]
  wire [26:0] _T_23; // @[RoundAnyRawFNToRecFN.scala 192:30:freechips.rocketchip.system.DefaultRV32Config.fir@190997.4]
  wire  _T_25; // @[RoundAnyRawFNToRecFN.scala 193:42:freechips.rocketchip.system.DefaultRV32Config.fir@190999.4]
  wire [25:0] _T_27; // @[RoundAnyRawFNToRecFN.scala 193:24:freechips.rocketchip.system.DefaultRV32Config.fir@191001.4]
  wire [25:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 192:47:freechips.rocketchip.system.DefaultRV32Config.fir@191002.4]
  wire [25:0] _T_28; // @[RoundAnyRawFNToRecFN.scala 192:47:freechips.rocketchip.system.DefaultRV32Config.fir@191002.4]
  wire [25:0] roundedSig; // @[RoundAnyRawFNToRecFN.scala 185:16:freechips.rocketchip.system.DefaultRV32Config.fir@191003.4]
  wire [2:0] _T_30; // @[RoundAnyRawFNToRecFN.scala 198:69:freechips.rocketchip.system.DefaultRV32Config.fir@191005.4]
  wire [9:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 198:40:freechips.rocketchip.system.DefaultRV32Config.fir@191006.4]
  wire [10:0] sRoundedExp; // @[RoundAnyRawFNToRecFN.scala 198:40:freechips.rocketchip.system.DefaultRV32Config.fir@191006.4]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 201:37:freechips.rocketchip.system.DefaultRV32Config.fir@191007.4]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 203:16:freechips.rocketchip.system.DefaultRV32Config.fir@191011.4]
  wire [3:0] _T_35; // @[RoundAnyRawFNToRecFN.scala 210:30:freechips.rocketchip.system.DefaultRV32Config.fir@191013.4]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 210:50:freechips.rocketchip.system.DefaultRV32Config.fir@191014.4]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 214:31:freechips.rocketchip.system.DefaultRV32Config.fir@191016.4]
  wire  unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 217:16:freechips.rocketchip.system.DefaultRV32Config.fir@191020.4]
  wire  _T_41; // @[RoundAnyRawFNToRecFN.scala 220:30:freechips.rocketchip.system.DefaultRV32Config.fir@191022.4]
  wire  _T_43; // @[RoundAnyRawFNToRecFN.scala 220:70:freechips.rocketchip.system.DefaultRV32Config.fir@191024.4]
  wire  unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 220:49:freechips.rocketchip.system.DefaultRV32Config.fir@191025.4]
  wire  _T_45; // @[RoundAnyRawFNToRecFN.scala 223:67:freechips.rocketchip.system.DefaultRV32Config.fir@191027.4]
  wire  _T_46; // @[RoundAnyRawFNToRecFN.scala 225:29:freechips.rocketchip.system.DefaultRV32Config.fir@191028.4]
  wire  unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 224:46:freechips.rocketchip.system.DefaultRV32Config.fir@191029.4]
  wire  roundCarry; // @[RoundAnyRawFNToRecFN.scala 228:16:freechips.rocketchip.system.DefaultRV32Config.fir@191032.4]
  wire [1:0] _T_49; // @[RoundAnyRawFNToRecFN.scala 238:48:freechips.rocketchip.system.DefaultRV32Config.fir@191033.4]
  wire  _T_50; // @[RoundAnyRawFNToRecFN.scala 238:62:freechips.rocketchip.system.DefaultRV32Config.fir@191034.4]
  wire  _T_51; // @[RoundAnyRawFNToRecFN.scala 238:32:freechips.rocketchip.system.DefaultRV32Config.fir@191035.4]
  wire  _T_54; // @[RoundAnyRawFNToRecFN.scala 239:30:freechips.rocketchip.system.DefaultRV32Config.fir@191038.4]
  wire  _T_55; // @[RoundAnyRawFNToRecFN.scala 238:74:freechips.rocketchip.system.DefaultRV32Config.fir@191039.4]
  wire  _T_59; // @[RoundAnyRawFNToRecFN.scala 241:39:freechips.rocketchip.system.DefaultRV32Config.fir@191043.4]
  wire  _T_60; // @[RoundAnyRawFNToRecFN.scala 241:34:freechips.rocketchip.system.DefaultRV32Config.fir@191044.4]
  wire  _T_62; // @[RoundAnyRawFNToRecFN.scala 244:38:freechips.rocketchip.system.DefaultRV32Config.fir@191046.4]
  wire  _T_63; // @[RoundAnyRawFNToRecFN.scala 245:45:freechips.rocketchip.system.DefaultRV32Config.fir@191047.4]
  wire  _T_64; // @[RoundAnyRawFNToRecFN.scala 245:60:freechips.rocketchip.system.DefaultRV32Config.fir@191048.4]
  wire  _T_65; // @[RoundAnyRawFNToRecFN.scala 240:27:freechips.rocketchip.system.DefaultRV32Config.fir@191049.4]
  wire  _T_66; // @[RoundAnyRawFNToRecFN.scala 239:76:freechips.rocketchip.system.DefaultRV32Config.fir@191050.4]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 235:40:freechips.rocketchip.system.DefaultRV32Config.fir@191051.4]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 248:49:freechips.rocketchip.system.DefaultRV32Config.fir@191053.4]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 253:34:freechips.rocketchip.system.DefaultRV32Config.fir@191055.4]
  wire  notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 254:49:freechips.rocketchip.system.DefaultRV32Config.fir@191056.4]
  wire  _T_69; // @[RoundAnyRawFNToRecFN.scala 255:22:freechips.rocketchip.system.DefaultRV32Config.fir@191057.4]
  wire  _T_70; // @[RoundAnyRawFNToRecFN.scala 255:36:freechips.rocketchip.system.DefaultRV32Config.fir@191058.4]
  wire  _T_71; // @[RoundAnyRawFNToRecFN.scala 255:33:freechips.rocketchip.system.DefaultRV32Config.fir@191059.4]
  wire  _T_72; // @[RoundAnyRawFNToRecFN.scala 255:64:freechips.rocketchip.system.DefaultRV32Config.fir@191060.4]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 255:61:freechips.rocketchip.system.DefaultRV32Config.fir@191061.4]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 256:32:freechips.rocketchip.system.DefaultRV32Config.fir@191062.4]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 257:32:freechips.rocketchip.system.DefaultRV32Config.fir@191063.4]
  wire  _T_73; // @[RoundAnyRawFNToRecFN.scala 258:43:freechips.rocketchip.system.DefaultRV32Config.fir@191064.4]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 258:28:freechips.rocketchip.system.DefaultRV32Config.fir@191065.4]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 261:60:freechips.rocketchip.system.DefaultRV32Config.fir@191067.4]
  wire  _T_75; // @[RoundAnyRawFNToRecFN.scala 263:20:freechips.rocketchip.system.DefaultRV32Config.fir@191068.4]
  wire  _T_76; // @[RoundAnyRawFNToRecFN.scala 263:60:freechips.rocketchip.system.DefaultRV32Config.fir@191069.4]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 263:45:freechips.rocketchip.system.DefaultRV32Config.fir@191070.4]
  wire  _T_77; // @[RoundAnyRawFNToRecFN.scala 264:42:freechips.rocketchip.system.DefaultRV32Config.fir@191071.4]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 264:39:freechips.rocketchip.system.DefaultRV32Config.fir@191072.4]
  wire  _T_78; // @[RoundAnyRawFNToRecFN.scala 266:45:freechips.rocketchip.system.DefaultRV32Config.fir@191073.4]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 266:32:freechips.rocketchip.system.DefaultRV32Config.fir@191074.4]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 268:22:freechips.rocketchip.system.DefaultRV32Config.fir@191075.4]
  wire  _T_79; // @[RoundAnyRawFNToRecFN.scala 271:32:freechips.rocketchip.system.DefaultRV32Config.fir@191076.4]
  wire [8:0] _T_80; // @[RoundAnyRawFNToRecFN.scala 271:18:freechips.rocketchip.system.DefaultRV32Config.fir@191077.4]
  wire [8:0] _T_81; // @[RoundAnyRawFNToRecFN.scala 271:14:freechips.rocketchip.system.DefaultRV32Config.fir@191078.4]
  wire [8:0] _T_82; // @[RoundAnyRawFNToRecFN.scala 270:24:freechips.rocketchip.system.DefaultRV32Config.fir@191079.4]
  wire [8:0] _T_84; // @[RoundAnyRawFNToRecFN.scala 275:18:freechips.rocketchip.system.DefaultRV32Config.fir@191081.4]
  wire [8:0] _T_85; // @[RoundAnyRawFNToRecFN.scala 275:14:freechips.rocketchip.system.DefaultRV32Config.fir@191082.4]
  wire [8:0] _T_86; // @[RoundAnyRawFNToRecFN.scala 274:17:freechips.rocketchip.system.DefaultRV32Config.fir@191083.4]
  wire [8:0] _T_87; // @[RoundAnyRawFNToRecFN.scala 279:18:freechips.rocketchip.system.DefaultRV32Config.fir@191084.4]
  wire [8:0] _T_88; // @[RoundAnyRawFNToRecFN.scala 279:14:freechips.rocketchip.system.DefaultRV32Config.fir@191085.4]
  wire [8:0] _T_89; // @[RoundAnyRawFNToRecFN.scala 278:17:freechips.rocketchip.system.DefaultRV32Config.fir@191086.4]
  wire [8:0] _T_90; // @[RoundAnyRawFNToRecFN.scala 283:18:freechips.rocketchip.system.DefaultRV32Config.fir@191087.4]
  wire [8:0] _T_91; // @[RoundAnyRawFNToRecFN.scala 283:14:freechips.rocketchip.system.DefaultRV32Config.fir@191088.4]
  wire [8:0] _T_92; // @[RoundAnyRawFNToRecFN.scala 282:17:freechips.rocketchip.system.DefaultRV32Config.fir@191089.4]
  wire [8:0] _T_93; // @[RoundAnyRawFNToRecFN.scala 287:16:freechips.rocketchip.system.DefaultRV32Config.fir@191090.4]
  wire [8:0] _T_94; // @[RoundAnyRawFNToRecFN.scala 286:18:freechips.rocketchip.system.DefaultRV32Config.fir@191091.4]
  wire [8:0] _T_95; // @[RoundAnyRawFNToRecFN.scala 291:16:freechips.rocketchip.system.DefaultRV32Config.fir@191092.4]
  wire [8:0] _T_96; // @[RoundAnyRawFNToRecFN.scala 290:15:freechips.rocketchip.system.DefaultRV32Config.fir@191093.4]
  wire [8:0] _T_97; // @[RoundAnyRawFNToRecFN.scala 295:16:freechips.rocketchip.system.DefaultRV32Config.fir@191094.4]
  wire [8:0] _T_98; // @[RoundAnyRawFNToRecFN.scala 294:15:freechips.rocketchip.system.DefaultRV32Config.fir@191095.4]
  wire [8:0] _T_99; // @[RoundAnyRawFNToRecFN.scala 296:16:freechips.rocketchip.system.DefaultRV32Config.fir@191096.4]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 295:77:freechips.rocketchip.system.DefaultRV32Config.fir@191097.4]
  wire  _T_100; // @[RoundAnyRawFNToRecFN.scala 298:22:freechips.rocketchip.system.DefaultRV32Config.fir@191098.4]
  wire  _T_101; // @[RoundAnyRawFNToRecFN.scala 298:38:freechips.rocketchip.system.DefaultRV32Config.fir@191099.4]
  wire [22:0] _T_102; // @[RoundAnyRawFNToRecFN.scala 299:16:freechips.rocketchip.system.DefaultRV32Config.fir@191100.4]
  wire [22:0] _T_103; // @[RoundAnyRawFNToRecFN.scala 298:12:freechips.rocketchip.system.DefaultRV32Config.fir@191101.4]
  wire [22:0] _T_105; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@191103.4]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 301:11:freechips.rocketchip.system.DefaultRV32Config.fir@191104.4]
  wire [9:0] _T_106; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@191105.4]
  wire [1:0] _T_108; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@191108.4]
  wire [2:0] _T_110; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@191110.4]
  my_lowMask my_lowMask ( // @[RoundAnyRawFNToRecFN.scala 160:40:freechips.rocketchip.system.DefaultRV32Config.fir@190967.4]
    .io_in(my_lowMask_io_in),
    .io_out(my_lowMask_io_out)
  );
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53:freechips.rocketchip.system.DefaultRV32Config.fir@190943.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53:freechips.rocketchip.system.DefaultRV32Config.fir@190945.4]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53:freechips.rocketchip.system.DefaultRV32Config.fir@190946.4]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53:freechips.rocketchip.system.DefaultRV32Config.fir@190947.4]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53:freechips.rocketchip.system.DefaultRV32Config.fir@190948.4]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27:freechips.rocketchip.system.DefaultRV32Config.fir@190949.4]
  assign _T_1 = ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:66:freechips.rocketchip.system.DefaultRV32Config.fir@190950.4]
  assign _T_2 = roundingMode_max & _T_1; // @[RoundAnyRawFNToRecFN.scala 96:63:freechips.rocketchip.system.DefaultRV32Config.fir@190951.4]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42:freechips.rocketchip.system.DefaultRV32Config.fir@190952.4]
  assign doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 120:61:freechips.rocketchip.system.DefaultRV32Config.fir@190954.4]
  assign _GEN_0 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 163:21:freechips.rocketchip.system.DefaultRV32Config.fir@190971.4]
  assign _T_4 = my_lowMask_io_out | _GEN_0; // @[RoundAnyRawFNToRecFN.scala 163:21:freechips.rocketchip.system.DefaultRV32Config.fir@190971.4]
  assign roundMask = {_T_4,2'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190972.4]
  assign shiftedRoundMask = {1'h0,roundMask[26:1]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190974.4]
  assign _T_6 = ~shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 170:28:freechips.rocketchip.system.DefaultRV32Config.fir@190975.4]
  assign roundPosMask = _T_6 & roundMask; // @[RoundAnyRawFNToRecFN.scala 170:46:freechips.rocketchip.system.DefaultRV32Config.fir@190976.4]
  assign _T_7 = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 172:40:freechips.rocketchip.system.DefaultRV32Config.fir@190977.4]
  assign roundPosBit = _T_7 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 172:56:freechips.rocketchip.system.DefaultRV32Config.fir@190978.4]
  assign _T_8 = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 174:42:freechips.rocketchip.system.DefaultRV32Config.fir@190979.4]
  assign anyRoundExtra = _T_8 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 174:62:freechips.rocketchip.system.DefaultRV32Config.fir@190980.4]
  assign anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 176:36:freechips.rocketchip.system.DefaultRV32Config.fir@190981.4]
  assign _T_9 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 180:38:freechips.rocketchip.system.DefaultRV32Config.fir@190982.4]
  assign _T_10 = _T_9 & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 180:67:freechips.rocketchip.system.DefaultRV32Config.fir@190983.4]
  assign _T_11 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 182:29:freechips.rocketchip.system.DefaultRV32Config.fir@190984.4]
  assign roundIncr = _T_10 | _T_11; // @[RoundAnyRawFNToRecFN.scala 181:31:freechips.rocketchip.system.DefaultRV32Config.fir@190985.4]
  assign _T_12 = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 186:32:freechips.rocketchip.system.DefaultRV32Config.fir@190986.4]
  assign _T_14 = _T_12[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 186:49:freechips.rocketchip.system.DefaultRV32Config.fir@190988.4]
  assign _T_15 = roundingMode_near_even & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 187:49:freechips.rocketchip.system.DefaultRV32Config.fir@190989.4]
  assign _T_16 = ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 188:30:freechips.rocketchip.system.DefaultRV32Config.fir@190990.4]
  assign _T_17 = _T_15 & _T_16; // @[RoundAnyRawFNToRecFN.scala 187:64:freechips.rocketchip.system.DefaultRV32Config.fir@190991.4]
  assign _T_19 = _T_17 ? roundMask[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 187:25:freechips.rocketchip.system.DefaultRV32Config.fir@190993.4]
  assign _T_20 = ~_T_19; // @[RoundAnyRawFNToRecFN.scala 187:21:freechips.rocketchip.system.DefaultRV32Config.fir@190994.4]
  assign _T_21 = _T_14 & _T_20; // @[RoundAnyRawFNToRecFN.scala 186:61:freechips.rocketchip.system.DefaultRV32Config.fir@190995.4]
  assign _T_22 = ~roundMask; // @[RoundAnyRawFNToRecFN.scala 192:32:freechips.rocketchip.system.DefaultRV32Config.fir@190996.4]
  assign _T_23 = io_in_sig & _T_22; // @[RoundAnyRawFNToRecFN.scala 192:30:freechips.rocketchip.system.DefaultRV32Config.fir@190997.4]
  assign _T_25 = roundingMode_odd & anyRound; // @[RoundAnyRawFNToRecFN.scala 193:42:freechips.rocketchip.system.DefaultRV32Config.fir@190999.4]
  assign _T_27 = _T_25 ? roundPosMask[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 193:24:freechips.rocketchip.system.DefaultRV32Config.fir@191001.4]
  assign _GEN_1 = {{1'd0}, _T_23[26:2]}; // @[RoundAnyRawFNToRecFN.scala 192:47:freechips.rocketchip.system.DefaultRV32Config.fir@191002.4]
  assign _T_28 = _GEN_1 | _T_27; // @[RoundAnyRawFNToRecFN.scala 192:47:freechips.rocketchip.system.DefaultRV32Config.fir@191002.4]
  assign roundedSig = roundIncr ? _T_21 : _T_28; // @[RoundAnyRawFNToRecFN.scala 185:16:freechips.rocketchip.system.DefaultRV32Config.fir@191003.4]
  assign _T_30 = {1'b0,$signed(roundedSig[25:24])}; // @[RoundAnyRawFNToRecFN.scala 198:69:freechips.rocketchip.system.DefaultRV32Config.fir@191005.4]
  assign _GEN_2 = {{7{_T_30[2]}},_T_30}; // @[RoundAnyRawFNToRecFN.scala 198:40:freechips.rocketchip.system.DefaultRV32Config.fir@191006.4]
  assign sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_2); // @[RoundAnyRawFNToRecFN.scala 198:40:freechips.rocketchip.system.DefaultRV32Config.fir@191006.4]
  assign common_expOut = sRoundedExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 201:37:freechips.rocketchip.system.DefaultRV32Config.fir@191007.4]
  assign common_fractOut = doShiftSigDown1 ? roundedSig[23:1] : roundedSig[22:0]; // @[RoundAnyRawFNToRecFN.scala 203:16:freechips.rocketchip.system.DefaultRV32Config.fir@191011.4]
  assign _T_35 = sRoundedExp[10:7]; // @[RoundAnyRawFNToRecFN.scala 210:30:freechips.rocketchip.system.DefaultRV32Config.fir@191013.4]
  assign common_overflow = $signed(_T_35) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 210:50:freechips.rocketchip.system.DefaultRV32Config.fir@191014.4]
  assign common_totalUnderflow = $signed(sRoundedExp) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 214:31:freechips.rocketchip.system.DefaultRV32Config.fir@191016.4]
  assign unboundedRange_roundPosBit = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 217:16:freechips.rocketchip.system.DefaultRV32Config.fir@191020.4]
  assign _T_41 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 220:30:freechips.rocketchip.system.DefaultRV32Config.fir@191022.4]
  assign _T_43 = io_in_sig[1:0] != 2'h0; // @[RoundAnyRawFNToRecFN.scala 220:70:freechips.rocketchip.system.DefaultRV32Config.fir@191024.4]
  assign unboundedRange_anyRound = _T_41 | _T_43; // @[RoundAnyRawFNToRecFN.scala 220:49:freechips.rocketchip.system.DefaultRV32Config.fir@191025.4]
  assign _T_45 = _T_9 & unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 223:67:freechips.rocketchip.system.DefaultRV32Config.fir@191027.4]
  assign _T_46 = roundMagUp & unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 225:29:freechips.rocketchip.system.DefaultRV32Config.fir@191028.4]
  assign unboundedRange_roundIncr = _T_45 | _T_46; // @[RoundAnyRawFNToRecFN.scala 224:46:freechips.rocketchip.system.DefaultRV32Config.fir@191029.4]
  assign roundCarry = doShiftSigDown1 ? roundedSig[25] : roundedSig[24]; // @[RoundAnyRawFNToRecFN.scala 228:16:freechips.rocketchip.system.DefaultRV32Config.fir@191032.4]
  assign _T_49 = io_in_sExp[9:8]; // @[RoundAnyRawFNToRecFN.scala 238:48:freechips.rocketchip.system.DefaultRV32Config.fir@191033.4]
  assign _T_50 = $signed(_T_49) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 238:62:freechips.rocketchip.system.DefaultRV32Config.fir@191034.4]
  assign _T_51 = anyRound & _T_50; // @[RoundAnyRawFNToRecFN.scala 238:32:freechips.rocketchip.system.DefaultRV32Config.fir@191035.4]
  assign _T_54 = doShiftSigDown1 ? roundMask[3] : roundMask[2]; // @[RoundAnyRawFNToRecFN.scala 239:30:freechips.rocketchip.system.DefaultRV32Config.fir@191038.4]
  assign _T_55 = _T_51 & _T_54; // @[RoundAnyRawFNToRecFN.scala 238:74:freechips.rocketchip.system.DefaultRV32Config.fir@191039.4]
  assign _T_59 = doShiftSigDown1 ? roundMask[4] : roundMask[3]; // @[RoundAnyRawFNToRecFN.scala 241:39:freechips.rocketchip.system.DefaultRV32Config.fir@191043.4]
  assign _T_60 = ~_T_59; // @[RoundAnyRawFNToRecFN.scala 241:34:freechips.rocketchip.system.DefaultRV32Config.fir@191044.4]
  assign _T_62 = _T_60 & roundCarry; // @[RoundAnyRawFNToRecFN.scala 244:38:freechips.rocketchip.system.DefaultRV32Config.fir@191046.4]
  assign _T_63 = _T_62 & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 245:45:freechips.rocketchip.system.DefaultRV32Config.fir@191047.4]
  assign _T_64 = _T_63 & unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 245:60:freechips.rocketchip.system.DefaultRV32Config.fir@191048.4]
  assign _T_65 = ~_T_64; // @[RoundAnyRawFNToRecFN.scala 240:27:freechips.rocketchip.system.DefaultRV32Config.fir@191049.4]
  assign _T_66 = _T_55 & _T_65; // @[RoundAnyRawFNToRecFN.scala 239:76:freechips.rocketchip.system.DefaultRV32Config.fir@191050.4]
  assign common_underflow = common_totalUnderflow | _T_66; // @[RoundAnyRawFNToRecFN.scala 235:40:freechips.rocketchip.system.DefaultRV32Config.fir@191051.4]
  assign common_inexact = common_totalUnderflow | anyRound; // @[RoundAnyRawFNToRecFN.scala 248:49:freechips.rocketchip.system.DefaultRV32Config.fir@191053.4]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 253:34:freechips.rocketchip.system.DefaultRV32Config.fir@191055.4]
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 254:49:freechips.rocketchip.system.DefaultRV32Config.fir@191056.4]
  assign _T_69 = ~isNaNOut; // @[RoundAnyRawFNToRecFN.scala 255:22:freechips.rocketchip.system.DefaultRV32Config.fir@191057.4]
  assign _T_70 = ~notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 255:36:freechips.rocketchip.system.DefaultRV32Config.fir@191058.4]
  assign _T_71 = _T_69 & _T_70; // @[RoundAnyRawFNToRecFN.scala 255:33:freechips.rocketchip.system.DefaultRV32Config.fir@191059.4]
  assign _T_72 = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 255:64:freechips.rocketchip.system.DefaultRV32Config.fir@191060.4]
  assign commonCase = _T_71 & _T_72; // @[RoundAnyRawFNToRecFN.scala 255:61:freechips.rocketchip.system.DefaultRV32Config.fir@191061.4]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 256:32:freechips.rocketchip.system.DefaultRV32Config.fir@191062.4]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 257:32:freechips.rocketchip.system.DefaultRV32Config.fir@191063.4]
  assign _T_73 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 258:43:freechips.rocketchip.system.DefaultRV32Config.fir@191064.4]
  assign inexact = overflow | _T_73; // @[RoundAnyRawFNToRecFN.scala 258:28:freechips.rocketchip.system.DefaultRV32Config.fir@191065.4]
  assign overflow_roundMagUp = _T_9 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 261:60:freechips.rocketchip.system.DefaultRV32Config.fir@191067.4]
  assign _T_75 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 263:20:freechips.rocketchip.system.DefaultRV32Config.fir@191068.4]
  assign _T_76 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 263:60:freechips.rocketchip.system.DefaultRV32Config.fir@191069.4]
  assign pegMinNonzeroMagOut = _T_75 & _T_76; // @[RoundAnyRawFNToRecFN.scala 263:45:freechips.rocketchip.system.DefaultRV32Config.fir@191070.4]
  assign _T_77 = ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 264:42:freechips.rocketchip.system.DefaultRV32Config.fir@191071.4]
  assign pegMaxFiniteMagOut = overflow & _T_77; // @[RoundAnyRawFNToRecFN.scala 264:39:freechips.rocketchip.system.DefaultRV32Config.fir@191072.4]
  assign _T_78 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 266:45:freechips.rocketchip.system.DefaultRV32Config.fir@191073.4]
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | _T_78; // @[RoundAnyRawFNToRecFN.scala 266:32:freechips.rocketchip.system.DefaultRV32Config.fir@191074.4]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 268:22:freechips.rocketchip.system.DefaultRV32Config.fir@191075.4]
  assign _T_79 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 271:32:freechips.rocketchip.system.DefaultRV32Config.fir@191076.4]
  assign _T_80 = _T_79 ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:18:freechips.rocketchip.system.DefaultRV32Config.fir@191077.4]
  assign _T_81 = ~_T_80; // @[RoundAnyRawFNToRecFN.scala 271:14:freechips.rocketchip.system.DefaultRV32Config.fir@191078.4]
  assign _T_82 = common_expOut & _T_81; // @[RoundAnyRawFNToRecFN.scala 270:24:freechips.rocketchip.system.DefaultRV32Config.fir@191079.4]
  assign _T_84 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:18:freechips.rocketchip.system.DefaultRV32Config.fir@191081.4]
  assign _T_85 = ~_T_84; // @[RoundAnyRawFNToRecFN.scala 275:14:freechips.rocketchip.system.DefaultRV32Config.fir@191082.4]
  assign _T_86 = _T_82 & _T_85; // @[RoundAnyRawFNToRecFN.scala 274:17:freechips.rocketchip.system.DefaultRV32Config.fir@191083.4]
  assign _T_87 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 279:18:freechips.rocketchip.system.DefaultRV32Config.fir@191084.4]
  assign _T_88 = ~_T_87; // @[RoundAnyRawFNToRecFN.scala 279:14:freechips.rocketchip.system.DefaultRV32Config.fir@191085.4]
  assign _T_89 = _T_86 & _T_88; // @[RoundAnyRawFNToRecFN.scala 278:17:freechips.rocketchip.system.DefaultRV32Config.fir@191086.4]
  assign _T_90 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 283:18:freechips.rocketchip.system.DefaultRV32Config.fir@191087.4]
  assign _T_91 = ~_T_90; // @[RoundAnyRawFNToRecFN.scala 283:14:freechips.rocketchip.system.DefaultRV32Config.fir@191088.4]
  assign _T_92 = _T_89 & _T_91; // @[RoundAnyRawFNToRecFN.scala 282:17:freechips.rocketchip.system.DefaultRV32Config.fir@191089.4]
  assign _T_93 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 287:16:freechips.rocketchip.system.DefaultRV32Config.fir@191090.4]
  assign _T_94 = _T_92 | _T_93; // @[RoundAnyRawFNToRecFN.scala 286:18:freechips.rocketchip.system.DefaultRV32Config.fir@191091.4]
  assign _T_95 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 291:16:freechips.rocketchip.system.DefaultRV32Config.fir@191092.4]
  assign _T_96 = _T_94 | _T_95; // @[RoundAnyRawFNToRecFN.scala 290:15:freechips.rocketchip.system.DefaultRV32Config.fir@191093.4]
  assign _T_97 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 295:16:freechips.rocketchip.system.DefaultRV32Config.fir@191094.4]
  assign _T_98 = _T_96 | _T_97; // @[RoundAnyRawFNToRecFN.scala 294:15:freechips.rocketchip.system.DefaultRV32Config.fir@191095.4]
  assign _T_99 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 296:16:freechips.rocketchip.system.DefaultRV32Config.fir@191096.4]
  assign expOut = _T_98 | _T_99; // @[RoundAnyRawFNToRecFN.scala 295:77:freechips.rocketchip.system.DefaultRV32Config.fir@191097.4]
  assign _T_100 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 298:22:freechips.rocketchip.system.DefaultRV32Config.fir@191098.4]
  assign _T_101 = _T_100 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 298:38:freechips.rocketchip.system.DefaultRV32Config.fir@191099.4]
  assign _T_102 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 299:16:freechips.rocketchip.system.DefaultRV32Config.fir@191100.4]
  assign _T_103 = _T_101 ? _T_102 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 298:12:freechips.rocketchip.system.DefaultRV32Config.fir@191101.4]
  assign _T_105 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@191103.4]
  assign fractOut = _T_103 | _T_105; // @[RoundAnyRawFNToRecFN.scala 301:11:freechips.rocketchip.system.DefaultRV32Config.fir@191104.4]
  assign _T_106 = {signOut,expOut}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@191105.4]
  assign _T_108 = {underflow,inexact}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@191108.4]
  assign _T_110 = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@191110.4]
  assign io_out = {_T_106,fractOut}; // @[RoundAnyRawFNToRecFN.scala 304:12:freechips.rocketchip.system.DefaultRV32Config.fir@191107.4]
  assign io_exceptionFlags = {_T_110,_T_108}; // @[RoundAnyRawFNToRecFN.scala 305:23:freechips.rocketchip.system.DefaultRV32Config.fir@191112.4]
  assign my_lowMask_io_in = io_in_sExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 161:34:freechips.rocketchip.system.DefaultRV32Config.fir@190970.4]
endmodule

module my_lowMask( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190850.2]
  input  [8:0]  io_in, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190851.4]
  output [24:0] io_out // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190851.4]
);
  wire [8:0] _T; // @[primitives.scala 54:40:freechips.rocketchip.system.DefaultRV32Config.fir@190854.4]
  wire  msb; // @[primitives.scala 126:25:freechips.rocketchip.system.DefaultRV32Config.fir@190855.4]
  wire [7:0] lsbs; // @[primitives.scala 128:26:freechips.rocketchip.system.DefaultRV32Config.fir@190856.4]
  wire  msb_1; // @[primitives.scala 126:25:freechips.rocketchip.system.DefaultRV32Config.fir@190857.4]
  wire [6:0] lsbs_1; // @[primitives.scala 128:26:freechips.rocketchip.system.DefaultRV32Config.fir@190858.4]
  wire  msb_2; // @[primitives.scala 126:25:freechips.rocketchip.system.DefaultRV32Config.fir@190859.4]
  wire [5:0] lsbs_2; // @[primitives.scala 128:26:freechips.rocketchip.system.DefaultRV32Config.fir@190860.4]
  wire [64:0] _T_1; // @[primitives.scala 163:58:freechips.rocketchip.system.DefaultRV32Config.fir@190861.4]
  wire [15:0] _T_7; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190867.4]
  wire [15:0] _T_9; // @[Bitwise.scala 102:65:freechips.rocketchip.system.DefaultRV32Config.fir@190869.4]
  wire [15:0] _T_11; // @[Bitwise.scala 102:75:freechips.rocketchip.system.DefaultRV32Config.fir@190871.4]
  wire [15:0] _T_12; // @[Bitwise.scala 102:39:freechips.rocketchip.system.DefaultRV32Config.fir@190872.4]
  wire [15:0] _GEN_0; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190877.4]
  wire [15:0] _T_17; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190877.4]
  wire [15:0] _T_19; // @[Bitwise.scala 102:65:freechips.rocketchip.system.DefaultRV32Config.fir@190879.4]
  wire [15:0] _T_21; // @[Bitwise.scala 102:75:freechips.rocketchip.system.DefaultRV32Config.fir@190881.4]
  wire [15:0] _T_22; // @[Bitwise.scala 102:39:freechips.rocketchip.system.DefaultRV32Config.fir@190882.4]
  wire [15:0] _GEN_1; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190887.4]
  wire [15:0] _T_27; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190887.4]
  wire [15:0] _T_29; // @[Bitwise.scala 102:65:freechips.rocketchip.system.DefaultRV32Config.fir@190889.4]
  wire [15:0] _T_31; // @[Bitwise.scala 102:75:freechips.rocketchip.system.DefaultRV32Config.fir@190891.4]
  wire [15:0] _T_32; // @[Bitwise.scala 102:39:freechips.rocketchip.system.DefaultRV32Config.fir@190892.4]
  wire [15:0] _GEN_2; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190897.4]
  wire [15:0] _T_37; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190897.4]
  wire [15:0] _T_39; // @[Bitwise.scala 102:65:freechips.rocketchip.system.DefaultRV32Config.fir@190899.4]
  wire [15:0] _T_41; // @[Bitwise.scala 102:75:freechips.rocketchip.system.DefaultRV32Config.fir@190901.4]
  wire [15:0] _T_42; // @[Bitwise.scala 102:39:freechips.rocketchip.system.DefaultRV32Config.fir@190902.4]
  wire [21:0] my_lowMask_1; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190919.4]
  wire [21:0] _T_59; // @[primitives.scala 159:25:freechips.rocketchip.system.DefaultRV32Config.fir@190920.4]
  wire [21:0] _T_60; // @[primitives.scala 157:21:freechips.rocketchip.system.DefaultRV32Config.fir@190921.4]
  wire [21:0] my_lowMask_1_1; // @[primitives.scala 157:17:freechips.rocketchip.system.DefaultRV32Config.fir@190922.4]
  wire [2:0] my_lowMask_1_2; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190932.4]
  wire [2:0] my_lowMask_2; // @[primitives.scala 134:24:freechips.rocketchip.system.DefaultRV32Config.fir@190933.4]
  wire [24:0] _T_68; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190934.4]
  wire [24:0] my_lowMask_1_3; // @[primitives.scala 144:24:freechips.rocketchip.system.DefaultRV32Config.fir@190935.4]
  assign _T = ~io_in; // @[primitives.scala 54:40:freechips.rocketchip.system.DefaultRV32Config.fir@190854.4]
  assign msb = _T[8]; // @[primitives.scala 126:25:freechips.rocketchip.system.DefaultRV32Config.fir@190855.4]
  assign lsbs = _T[7:0]; // @[primitives.scala 128:26:freechips.rocketchip.system.DefaultRV32Config.fir@190856.4]
  assign msb_1 = lsbs[7]; // @[primitives.scala 126:25:freechips.rocketchip.system.DefaultRV32Config.fir@190857.4]
  assign lsbs_1 = lsbs[6:0]; // @[primitives.scala 128:26:freechips.rocketchip.system.DefaultRV32Config.fir@190858.4]
  assign msb_2 = lsbs_1[6]; // @[primitives.scala 126:25:freechips.rocketchip.system.DefaultRV32Config.fir@190859.4]
  assign lsbs_2 = lsbs_1[5:0]; // @[primitives.scala 128:26:freechips.rocketchip.system.DefaultRV32Config.fir@190860.4]
  assign _T_1 = -65'sh10000000000000000 >>> lsbs_2; // @[primitives.scala 163:58:freechips.rocketchip.system.DefaultRV32Config.fir@190861.4]
  assign _T_7 = {{8'd0}, _T_1[57:50]}; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190867.4]
  assign _T_9 = {_T_1[49:42], 8'h0}; // @[Bitwise.scala 102:65:freechips.rocketchip.system.DefaultRV32Config.fir@190869.4]
  assign _T_11 = _T_9 & 16'hff00; // @[Bitwise.scala 102:75:freechips.rocketchip.system.DefaultRV32Config.fir@190871.4]
  assign _T_12 = _T_7 | _T_11; // @[Bitwise.scala 102:39:freechips.rocketchip.system.DefaultRV32Config.fir@190872.4]
  assign _GEN_0 = {{4'd0}, _T_12[15:4]}; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190877.4]
  assign _T_17 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190877.4]
  assign _T_19 = {_T_12[11:0], 4'h0}; // @[Bitwise.scala 102:65:freechips.rocketchip.system.DefaultRV32Config.fir@190879.4]
  assign _T_21 = _T_19 & 16'hf0f0; // @[Bitwise.scala 102:75:freechips.rocketchip.system.DefaultRV32Config.fir@190881.4]
  assign _T_22 = _T_17 | _T_21; // @[Bitwise.scala 102:39:freechips.rocketchip.system.DefaultRV32Config.fir@190882.4]
  assign _GEN_1 = {{2'd0}, _T_22[15:2]}; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190887.4]
  assign _T_27 = _GEN_1 & 16'h3333; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190887.4]
  assign _T_29 = {_T_22[13:0], 2'h0}; // @[Bitwise.scala 102:65:freechips.rocketchip.system.DefaultRV32Config.fir@190889.4]
  assign _T_31 = _T_29 & 16'hcccc; // @[Bitwise.scala 102:75:freechips.rocketchip.system.DefaultRV32Config.fir@190891.4]
  assign _T_32 = _T_27 | _T_31; // @[Bitwise.scala 102:39:freechips.rocketchip.system.DefaultRV32Config.fir@190892.4]
  assign _GEN_2 = {{1'd0}, _T_32[15:1]}; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190897.4]
  assign _T_37 = _GEN_2 & 16'h5555; // @[Bitwise.scala 102:31:freechips.rocketchip.system.DefaultRV32Config.fir@190897.4]
  assign _T_39 = {_T_32[14:0], 1'h0}; // @[Bitwise.scala 102:65:freechips.rocketchip.system.DefaultRV32Config.fir@190899.4]
  assign _T_41 = _T_39 & 16'haaaa; // @[Bitwise.scala 102:75:freechips.rocketchip.system.DefaultRV32Config.fir@190901.4]
  assign _T_42 = _T_37 | _T_41; // @[Bitwise.scala 102:39:freechips.rocketchip.system.DefaultRV32Config.fir@190902.4]
  assign my_lowMask_1 = {_T_42,_T_1[58],_T_1[59],_T_1[60],_T_1[61],_T_1[62],_T_1[63]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190919.4]
  assign _T_59 = ~my_lowMask_1; // @[primitives.scala 159:25:freechips.rocketchip.system.DefaultRV32Config.fir@190920.4]
  assign _T_60 = msb_2 ? 22'h0 : _T_59; // @[primitives.scala 157:21:freechips.rocketchip.system.DefaultRV32Config.fir@190921.4]
  assign my_lowMask_1_1 = ~_T_60; // @[primitives.scala 157:17:freechips.rocketchip.system.DefaultRV32Config.fir@190922.4]
  assign my_lowMask_1_2 = {_T_1[0],_T_1[1],_T_1[2]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190932.4]
  assign my_lowMask_2 = msb_2 ? my_lowMask_1_2 : 3'h0; // @[primitives.scala 134:24:freechips.rocketchip.system.DefaultRV32Config.fir@190933.4]
  assign _T_68 = {my_lowMask_1_1,3'h7}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190934.4]
  assign my_lowMask_1_3 = msb_1 ? _T_68 : {{22'd0}, my_lowMask_2}; // @[primitives.scala 144:24:freechips.rocketchip.system.DefaultRV32Config.fir@190935.4]
  assign io_out = msb ? my_lowMask_1_3 : 25'h0; // @[primitives.scala 106:16:freechips.rocketchip.system.DefaultRV32Config.fir@190937.4]
endmodule

