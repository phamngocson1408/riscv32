module MulAddRecFNToRaw_preMul( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190274.2]
  input  [1:0]  io_op, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  input  [32:0] io_a, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  input  [32:0] io_b, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  input  [32:0] io_c, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output [23:0] io_mulAddA, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output [23:0] io_mulAddB, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output [47:0] io_mulAddC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isSigNaNAny, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isNaNAOrB, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isInfA, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isZeroA, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isInfB, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isZeroB, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_signProd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isNaNC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isInfC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_isZeroC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output [9:0]  io_toPostMul_sExpSum, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_doSubMags, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_CIsDominant, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output [4:0]  io_toPostMul_CDom_CAlignDist, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output [25:0] io_toPostMul_highAlignedSigC, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
  output        io_toPostMul_bit0AlignedSigC // @[:freechips.rocketchip.system.DefaultRV32Config.fir@190275.4]
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@190280.4]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@190282.4]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@190286.4]
  wire  _T_8; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@190289.4]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@190293.4]
  wire [9:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@190295.4]
  wire  _T_12; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@190297.4]
  wire [24:0] rawA_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190300.4]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@190304.4]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@190306.4]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@190310.4]
  wire  _T_24; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@190313.4]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@190317.4]
  wire [9:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@190319.4]
  wire  _T_28; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@190321.4]
  wire [24:0] rawB_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190324.4]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@190328.4]
  wire  _T_36; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@190330.4]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@190334.4]
  wire  _T_40; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@190337.4]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@190341.4]
  wire [9:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@190343.4]
  wire  _T_44; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@190345.4]
  wire [24:0] rawC_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190348.4]
  wire  _T_48; // @[MulAddRecFN.scala 98:30:freechips.rocketchip.system.DefaultRV32Config.fir@190350.4]
  wire  signProd; // @[MulAddRecFN.scala 98:42:freechips.rocketchip.system.DefaultRV32Config.fir@190352.4]
  wire [10:0] _T_50; // @[MulAddRecFN.scala 101:19:freechips.rocketchip.system.DefaultRV32Config.fir@190353.4]
  wire [10:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32:freechips.rocketchip.system.DefaultRV32Config.fir@190356.4]
  wire  _T_53; // @[MulAddRecFN.scala 103:30:freechips.rocketchip.system.DefaultRV32Config.fir@190357.4]
  wire  doSubMags; // @[MulAddRecFN.scala 103:42:freechips.rocketchip.system.DefaultRV32Config.fir@190359.4]
  wire [10:0] _GEN_0; // @[MulAddRecFN.scala 107:42:freechips.rocketchip.system.DefaultRV32Config.fir@190360.4]
  wire [10:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42:freechips.rocketchip.system.DefaultRV32Config.fir@190362.4]
  wire [9:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42:freechips.rocketchip.system.DefaultRV32Config.fir@190363.4]
  wire  _T_57; // @[MulAddRecFN.scala 109:35:freechips.rocketchip.system.DefaultRV32Config.fir@190364.4]
  wire  _T_58; // @[MulAddRecFN.scala 109:69:freechips.rocketchip.system.DefaultRV32Config.fir@190365.4]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50:freechips.rocketchip.system.DefaultRV32Config.fir@190366.4]
  wire  _T_60; // @[MulAddRecFN.scala 111:60:freechips.rocketchip.system.DefaultRV32Config.fir@190368.4]
  wire  _T_61; // @[MulAddRecFN.scala 111:39:freechips.rocketchip.system.DefaultRV32Config.fir@190369.4]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23:freechips.rocketchip.system.DefaultRV32Config.fir@190370.4]
  wire  _T_62; // @[MulAddRecFN.scala 115:34:freechips.rocketchip.system.DefaultRV32Config.fir@190371.4]
  wire [6:0] _T_64; // @[MulAddRecFN.scala 115:16:freechips.rocketchip.system.DefaultRV32Config.fir@190373.4]
  wire [6:0] CAlignDist; // @[MulAddRecFN.scala 113:12:freechips.rocketchip.system.DefaultRV32Config.fir@190374.4]
  wire [24:0] _T_65; // @[MulAddRecFN.scala 121:28:freechips.rocketchip.system.DefaultRV32Config.fir@190375.4]
  wire [24:0] _T_66; // @[MulAddRecFN.scala 121:16:freechips.rocketchip.system.DefaultRV32Config.fir@190376.4]
  wire [52:0] _T_68; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@190378.4]
  wire [77:0] _T_70; // @[MulAddRecFN.scala 123:11:freechips.rocketchip.system.DefaultRV32Config.fir@190380.4]
  wire [77:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17:freechips.rocketchip.system.DefaultRV32Config.fir@190381.4]
  wire [26:0] _T_71; // @[MulAddRecFN.scala 125:30:freechips.rocketchip.system.DefaultRV32Config.fir@190382.4]
  wire  _T_74; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190386.4]
  wire  _T_76; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190389.4]
  wire  _T_78; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190392.4]
  wire  _T_80; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190395.4]
  wire  _T_82; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190398.4]
  wire  _T_84; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190401.4]
  wire  _T_86; // @[primitives.scala 208:57:freechips.rocketchip.system.DefaultRV32Config.fir@190404.4]
  wire [6:0] _T_92; // @[primitives.scala 209:20:freechips.rocketchip.system.DefaultRV32Config.fir@190411.4]
  wire [32:0] shift; // @[primitives.scala 160:58:freechips.rocketchip.system.DefaultRV32Config.fir@190413.4]
  wire [5:0] _T_109; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190429.4]
  wire [6:0] _GEN_1; // @[MulAddRecFN.scala 125:68:freechips.rocketchip.system.DefaultRV32Config.fir@190430.4]
  wire [6:0] _T_110; // @[MulAddRecFN.scala 125:68:freechips.rocketchip.system.DefaultRV32Config.fir@190430.4]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11:freechips.rocketchip.system.DefaultRV32Config.fir@190431.4]
  wire  _T_113; // @[MulAddRecFN.scala 137:39:freechips.rocketchip.system.DefaultRV32Config.fir@190434.4]
  wire  _T_114; // @[MulAddRecFN.scala 137:47:freechips.rocketchip.system.DefaultRV32Config.fir@190435.4]
  wire  _T_115; // @[MulAddRecFN.scala 137:44:freechips.rocketchip.system.DefaultRV32Config.fir@190436.4]
  wire  _T_117; // @[MulAddRecFN.scala 138:39:freechips.rocketchip.system.DefaultRV32Config.fir@190438.4]
  wire  _T_118; // @[MulAddRecFN.scala 138:44:freechips.rocketchip.system.DefaultRV32Config.fir@190439.4]
  wire  _T_119; // @[MulAddRecFN.scala 136:16:freechips.rocketchip.system.DefaultRV32Config.fir@190440.4]
  wire [74:0] _T_120; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190441.4]
  wire [75:0] alignedSigC; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190442.4]
  wire  _T_123; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@190448.4]
  wire  _T_124; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@190449.4]
  wire  _T_126; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@190451.4]
  wire  _T_127; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@190452.4]
  wire  _T_128; // @[MulAddRecFN.scala 149:32:freechips.rocketchip.system.DefaultRV32Config.fir@190453.4]
  wire  _T_130; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@190455.4]
  wire  _T_131; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@190456.4]
  wire [10:0] _T_136; // @[MulAddRecFN.scala 161:53:freechips.rocketchip.system.DefaultRV32Config.fir@190471.4]
  wire [10:0] _T_137; // @[MulAddRecFN.scala 161:12:freechips.rocketchip.system.DefaultRV32Config.fir@190472.4]
  assign rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@190280.4]
  assign _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@190282.4]
  assign rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@190286.4]
  assign _T_8 = ~io_a[29]; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@190289.4]
  assign rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@190293.4]
  assign rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@190295.4]
  assign _T_12 = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@190297.4]
  assign rawA_sig = {1'h0,_T_12,io_a[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190300.4]
  assign rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@190304.4]
  assign _T_20 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@190306.4]
  assign rawB_isNaN = _T_20 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@190310.4]
  assign _T_24 = ~io_b[29]; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@190313.4]
  assign rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@190317.4]
  assign rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@190319.4]
  assign _T_28 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@190321.4]
  assign rawB_sig = {1'h0,_T_28,io_b[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190324.4]
  assign rawC_isZero = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@190328.4]
  assign _T_36 = io_c[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@190330.4]
  assign rawC_isNaN = _T_36 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@190334.4]
  assign _T_40 = ~io_c[29]; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@190337.4]
  assign rawC_sign = io_c[32]; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@190341.4]
  assign rawC_sExp = {1'b0,$signed(io_c[31:23])}; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@190343.4]
  assign _T_44 = ~rawC_isZero; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@190345.4]
  assign rawC_sig = {1'h0,_T_44,io_c[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190348.4]
  assign _T_48 = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30:freechips.rocketchip.system.DefaultRV32Config.fir@190350.4]
  assign signProd = _T_48 ^ io_op[1]; // @[MulAddRecFN.scala 98:42:freechips.rocketchip.system.DefaultRV32Config.fir@190352.4]
  assign _T_50 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19:freechips.rocketchip.system.DefaultRV32Config.fir@190353.4]
  assign sExpAlignedProd = $signed(_T_50) - 11'she5; // @[MulAddRecFN.scala 101:32:freechips.rocketchip.system.DefaultRV32Config.fir@190356.4]
  assign _T_53 = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30:freechips.rocketchip.system.DefaultRV32Config.fir@190357.4]
  assign doSubMags = _T_53 ^ io_op[0]; // @[MulAddRecFN.scala 103:42:freechips.rocketchip.system.DefaultRV32Config.fir@190359.4]
  assign _GEN_0 = {{1{rawC_sExp[9]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42:freechips.rocketchip.system.DefaultRV32Config.fir@190360.4]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42:freechips.rocketchip.system.DefaultRV32Config.fir@190362.4]
  assign posNatCAlignDist = sNatCAlignDist[9:0]; // @[MulAddRecFN.scala 108:42:freechips.rocketchip.system.DefaultRV32Config.fir@190363.4]
  assign _T_57 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35:freechips.rocketchip.system.DefaultRV32Config.fir@190364.4]
  assign _T_58 = $signed(sNatCAlignDist) < 11'sh0; // @[MulAddRecFN.scala 109:69:freechips.rocketchip.system.DefaultRV32Config.fir@190365.4]
  assign isMinCAlign = _T_57 | _T_58; // @[MulAddRecFN.scala 109:50:freechips.rocketchip.system.DefaultRV32Config.fir@190366.4]
  assign _T_60 = posNatCAlignDist <= 10'h18; // @[MulAddRecFN.scala 111:60:freechips.rocketchip.system.DefaultRV32Config.fir@190368.4]
  assign _T_61 = isMinCAlign | _T_60; // @[MulAddRecFN.scala 111:39:freechips.rocketchip.system.DefaultRV32Config.fir@190369.4]
  assign CIsDominant = _T_44 & _T_61; // @[MulAddRecFN.scala 111:23:freechips.rocketchip.system.DefaultRV32Config.fir@190370.4]
  assign _T_62 = posNatCAlignDist < 10'h4a; // @[MulAddRecFN.scala 115:34:freechips.rocketchip.system.DefaultRV32Config.fir@190371.4]
  assign _T_64 = _T_62 ? posNatCAlignDist[6:0] : 7'h4a; // @[MulAddRecFN.scala 115:16:freechips.rocketchip.system.DefaultRV32Config.fir@190373.4]
  assign CAlignDist = isMinCAlign ? 7'h0 : _T_64; // @[MulAddRecFN.scala 113:12:freechips.rocketchip.system.DefaultRV32Config.fir@190374.4]
  assign _T_65 = ~rawC_sig; // @[MulAddRecFN.scala 121:28:freechips.rocketchip.system.DefaultRV32Config.fir@190375.4]
  assign _T_66 = doSubMags ? _T_65 : rawC_sig; // @[MulAddRecFN.scala 121:16:freechips.rocketchip.system.DefaultRV32Config.fir@190376.4]
  assign _T_68 = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 71:12:freechips.rocketchip.system.DefaultRV32Config.fir@190378.4]
  assign _T_70 = {_T_66,_T_68}; // @[MulAddRecFN.scala 123:11:freechips.rocketchip.system.DefaultRV32Config.fir@190380.4]
  assign mainAlignedSigC = $signed(_T_70) >>> CAlignDist; // @[MulAddRecFN.scala 123:17:freechips.rocketchip.system.DefaultRV32Config.fir@190381.4]
  assign _T_71 = {rawC_sig, 2'h0}; // @[MulAddRecFN.scala 125:30:freechips.rocketchip.system.DefaultRV32Config.fir@190382.4]
  assign _T_74 = _T_71[3:0] != 4'h0; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190386.4]
  assign _T_76 = _T_71[7:4] != 4'h0; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190389.4]
  assign _T_78 = _T_71[11:8] != 4'h0; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190392.4]
  assign _T_80 = _T_71[15:12] != 4'h0; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190395.4]
  assign _T_82 = _T_71[19:16] != 4'h0; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190398.4]
  assign _T_84 = _T_71[23:20] != 4'h0; // @[primitives.scala 205:54:freechips.rocketchip.system.DefaultRV32Config.fir@190401.4]
  assign _T_86 = _T_71[26:24] != 3'h0; // @[primitives.scala 208:57:freechips.rocketchip.system.DefaultRV32Config.fir@190404.4]
  assign _T_92 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76,_T_74}; // @[primitives.scala 209:20:freechips.rocketchip.system.DefaultRV32Config.fir@190411.4]
  assign shift = -33'sh100000000 >>> CAlignDist[6:2]; // @[primitives.scala 160:58:freechips.rocketchip.system.DefaultRV32Config.fir@190413.4]
  assign _T_109 = {shift[14],shift[15],shift[16],shift[17],shift[18],shift[19]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190429.4]
  assign _GEN_1 = {{1'd0}, _T_109}; // @[MulAddRecFN.scala 125:68:freechips.rocketchip.system.DefaultRV32Config.fir@190430.4]
  assign _T_110 = _T_92 & _GEN_1; // @[MulAddRecFN.scala 125:68:freechips.rocketchip.system.DefaultRV32Config.fir@190430.4]
  assign reduced4CExtra = _T_110 != 7'h0; // @[MulAddRecFN.scala 133:11:freechips.rocketchip.system.DefaultRV32Config.fir@190431.4]
  assign _T_113 = mainAlignedSigC[2:0] == 3'h7; // @[MulAddRecFN.scala 137:39:freechips.rocketchip.system.DefaultRV32Config.fir@190434.4]
  assign _T_114 = ~reduced4CExtra; // @[MulAddRecFN.scala 137:47:freechips.rocketchip.system.DefaultRV32Config.fir@190435.4]
  assign _T_115 = _T_113 & _T_114; // @[MulAddRecFN.scala 137:44:freechips.rocketchip.system.DefaultRV32Config.fir@190436.4]
  assign _T_117 = mainAlignedSigC[2:0] != 3'h0; // @[MulAddRecFN.scala 138:39:freechips.rocketchip.system.DefaultRV32Config.fir@190438.4]
  assign _T_118 = _T_117 | reduced4CExtra; // @[MulAddRecFN.scala 138:44:freechips.rocketchip.system.DefaultRV32Config.fir@190439.4]
  assign _T_119 = doSubMags ? _T_115 : _T_118; // @[MulAddRecFN.scala 136:16:freechips.rocketchip.system.DefaultRV32Config.fir@190440.4]
  assign _T_120 = mainAlignedSigC[77:3]; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190441.4]
  assign alignedSigC = {_T_120,_T_119}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@190442.4]
  assign _T_123 = ~rawA_sig[22]; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@190448.4]
  assign _T_124 = rawA_isNaN & _T_123; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@190449.4]
  assign _T_126 = ~rawB_sig[22]; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@190451.4]
  assign _T_127 = rawB_isNaN & _T_126; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@190452.4]
  assign _T_128 = _T_124 | _T_127; // @[MulAddRecFN.scala 149:32:freechips.rocketchip.system.DefaultRV32Config.fir@190453.4]
  assign _T_130 = ~rawC_sig[22]; // @[common.scala 81:49:freechips.rocketchip.system.DefaultRV32Config.fir@190455.4]
  assign _T_131 = rawC_isNaN & _T_130; // @[common.scala 81:46:freechips.rocketchip.system.DefaultRV32Config.fir@190456.4]
  assign _T_136 = $signed(sExpAlignedProd) - 11'sh18; // @[MulAddRecFN.scala 161:53:freechips.rocketchip.system.DefaultRV32Config.fir@190471.4]
  assign _T_137 = CIsDominant ? $signed({{1{rawC_sExp[9]}},rawC_sExp}) : $signed(_T_136); // @[MulAddRecFN.scala 161:12:freechips.rocketchip.system.DefaultRV32Config.fir@190472.4]
  assign io_mulAddA = rawA_sig[23:0]; // @[MulAddRecFN.scala 144:16:freechips.rocketchip.system.DefaultRV32Config.fir@190443.4]
  assign io_mulAddB = rawB_sig[23:0]; // @[MulAddRecFN.scala 145:16:freechips.rocketchip.system.DefaultRV32Config.fir@190444.4]
  assign io_mulAddC = alignedSigC[48:1]; // @[MulAddRecFN.scala 146:16:freechips.rocketchip.system.DefaultRV32Config.fir@190446.4]
  assign io_toPostMul_isSigNaNAny = _T_128 | _T_131; // @[MulAddRecFN.scala 148:30:freechips.rocketchip.system.DefaultRV32Config.fir@190458.4]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28:freechips.rocketchip.system.DefaultRV32Config.fir@190460.4]
  assign io_toPostMul_isInfA = _T_4 & _T_8; // @[MulAddRecFN.scala 152:28:freechips.rocketchip.system.DefaultRV32Config.fir@190461.4]
  assign io_toPostMul_isZeroA = io_a[31:29] == 3'h0; // @[MulAddRecFN.scala 153:28:freechips.rocketchip.system.DefaultRV32Config.fir@190462.4]
  assign io_toPostMul_isInfB = _T_20 & _T_24; // @[MulAddRecFN.scala 154:28:freechips.rocketchip.system.DefaultRV32Config.fir@190463.4]
  assign io_toPostMul_isZeroB = io_b[31:29] == 3'h0; // @[MulAddRecFN.scala 155:28:freechips.rocketchip.system.DefaultRV32Config.fir@190464.4]
  assign io_toPostMul_signProd = _T_48 ^ io_op[1]; // @[MulAddRecFN.scala 156:28:freechips.rocketchip.system.DefaultRV32Config.fir@190465.4]
  assign io_toPostMul_isNaNC = _T_36 & io_c[29]; // @[MulAddRecFN.scala 157:28:freechips.rocketchip.system.DefaultRV32Config.fir@190466.4]
  assign io_toPostMul_isInfC = _T_36 & _T_40; // @[MulAddRecFN.scala 158:28:freechips.rocketchip.system.DefaultRV32Config.fir@190467.4]
  assign io_toPostMul_isZeroC = io_c[31:29] == 3'h0; // @[MulAddRecFN.scala 159:28:freechips.rocketchip.system.DefaultRV32Config.fir@190468.4]
  assign io_toPostMul_sExpSum = _T_137[9:0]; // @[MulAddRecFN.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@190473.4]
  assign io_toPostMul_doSubMags = _T_53 ^ io_op[0]; // @[MulAddRecFN.scala 162:28:freechips.rocketchip.system.DefaultRV32Config.fir@190474.4]
  assign io_toPostMul_CIsDominant = _T_44 & _T_61; // @[MulAddRecFN.scala 163:30:freechips.rocketchip.system.DefaultRV32Config.fir@190475.4]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[MulAddRecFN.scala 164:34:freechips.rocketchip.system.DefaultRV32Config.fir@190477.4]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[MulAddRecFN.scala 165:34:freechips.rocketchip.system.DefaultRV32Config.fir@190479.4]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34:freechips.rocketchip.system.DefaultRV32Config.fir@190481.4]
endmodule

