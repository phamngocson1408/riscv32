module RoundAnyRawFNToRecFN_1( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@173374.2]
  input         io_in_isZero, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@173375.4]
  input         io_in_sign, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@173375.4]
  input  [7:0]  io_in_sExp, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@173375.4]
  input  [32:0] io_in_sig, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@173375.4]
  input  [2:0]  io_roundingMode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@173375.4]
  output [32:0] io_out, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@173375.4]
  output [4:0]  io_exceptionFlags // @[:freechips.rocketchip.system.DefaultRV32Config.fir@173375.4]
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53:freechips.rocketchip.system.DefaultRV32Config.fir@173378.4]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53:freechips.rocketchip.system.DefaultRV32Config.fir@173380.4]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53:freechips.rocketchip.system.DefaultRV32Config.fir@173381.4]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53:freechips.rocketchip.system.DefaultRV32Config.fir@173382.4]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53:freechips.rocketchip.system.DefaultRV32Config.fir@173383.4]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27:freechips.rocketchip.system.DefaultRV32Config.fir@173384.4]
  wire  _T_1; // @[RoundAnyRawFNToRecFN.scala 96:66:freechips.rocketchip.system.DefaultRV32Config.fir@173385.4]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63:freechips.rocketchip.system.DefaultRV32Config.fir@173386.4]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42:freechips.rocketchip.system.DefaultRV32Config.fir@173387.4]
  wire [8:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@173388.4]
  wire [9:0] _T_3; // @[RoundAnyRawFNToRecFN.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@173388.4]
  wire [8:0] _T_4; // @[RoundAnyRawFNToRecFN.scala 104:14:freechips.rocketchip.system.DefaultRV32Config.fir@173389.4]
  wire [9:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31:freechips.rocketchip.system.DefaultRV32Config.fir@173390.4]
  wire [25:0] _T_5; // @[RoundAnyRawFNToRecFN.scala 115:26:freechips.rocketchip.system.DefaultRV32Config.fir@173391.4]
  wire [6:0] _T_6; // @[RoundAnyRawFNToRecFN.scala 116:26:freechips.rocketchip.system.DefaultRV32Config.fir@173392.4]
  wire  _T_7; // @[RoundAnyRawFNToRecFN.scala 116:60:freechips.rocketchip.system.DefaultRV32Config.fir@173393.4]
  wire [26:0] adjustedSig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@173394.4]
  wire [26:0] _T_11; // @[RoundAnyRawFNToRecFN.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@173413.4]
  wire  roundPosBit; // @[RoundAnyRawFNToRecFN.scala 173:56:freechips.rocketchip.system.DefaultRV32Config.fir@173414.4]
  wire [26:0] _T_12; // @[RoundAnyRawFNToRecFN.scala 175:42:freechips.rocketchip.system.DefaultRV32Config.fir@173415.4]
  wire  anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 175:62:freechips.rocketchip.system.DefaultRV32Config.fir@173416.4]
  wire  anyRound; // @[RoundAnyRawFNToRecFN.scala 177:36:freechips.rocketchip.system.DefaultRV32Config.fir@173417.4]
  wire  _T_13; // @[RoundAnyRawFNToRecFN.scala 181:38:freechips.rocketchip.system.DefaultRV32Config.fir@173418.4]
  wire  _T_14; // @[RoundAnyRawFNToRecFN.scala 181:67:freechips.rocketchip.system.DefaultRV32Config.fir@173419.4]
  wire  _T_15; // @[RoundAnyRawFNToRecFN.scala 183:29:freechips.rocketchip.system.DefaultRV32Config.fir@173420.4]
  wire  roundIncr; // @[RoundAnyRawFNToRecFN.scala 182:31:freechips.rocketchip.system.DefaultRV32Config.fir@173421.4]
  wire [26:0] _T_16; // @[RoundAnyRawFNToRecFN.scala 187:32:freechips.rocketchip.system.DefaultRV32Config.fir@173422.4]
  wire [24:0] _T_17; // @[RoundAnyRawFNToRecFN.scala 187:44:freechips.rocketchip.system.DefaultRV32Config.fir@173423.4]
  wire [25:0] _T_18; // @[RoundAnyRawFNToRecFN.scala 187:49:freechips.rocketchip.system.DefaultRV32Config.fir@173424.4]
  wire  _T_19; // @[RoundAnyRawFNToRecFN.scala 188:49:freechips.rocketchip.system.DefaultRV32Config.fir@173425.4]
  wire  _T_20; // @[RoundAnyRawFNToRecFN.scala 189:30:freechips.rocketchip.system.DefaultRV32Config.fir@173426.4]
  wire  _T_21; // @[RoundAnyRawFNToRecFN.scala 188:64:freechips.rocketchip.system.DefaultRV32Config.fir@173427.4]
  wire [25:0] _T_23; // @[RoundAnyRawFNToRecFN.scala 188:25:freechips.rocketchip.system.DefaultRV32Config.fir@173429.4]
  wire [25:0] _T_24; // @[RoundAnyRawFNToRecFN.scala 188:21:freechips.rocketchip.system.DefaultRV32Config.fir@173430.4]
  wire [25:0] _T_25; // @[RoundAnyRawFNToRecFN.scala 187:61:freechips.rocketchip.system.DefaultRV32Config.fir@173431.4]
  wire [26:0] _T_27; // @[RoundAnyRawFNToRecFN.scala 193:30:freechips.rocketchip.system.DefaultRV32Config.fir@173433.4]
  wire [24:0] _T_28; // @[RoundAnyRawFNToRecFN.scala 193:43:freechips.rocketchip.system.DefaultRV32Config.fir@173434.4]
  wire  _T_29; // @[RoundAnyRawFNToRecFN.scala 194:42:freechips.rocketchip.system.DefaultRV32Config.fir@173435.4]
  wire [25:0] _T_31; // @[RoundAnyRawFNToRecFN.scala 194:24:freechips.rocketchip.system.DefaultRV32Config.fir@173437.4]
  wire [25:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 193:47:freechips.rocketchip.system.DefaultRV32Config.fir@173438.4]
  wire [25:0] _T_32; // @[RoundAnyRawFNToRecFN.scala 193:47:freechips.rocketchip.system.DefaultRV32Config.fir@173438.4]
  wire [25:0] roundedSig; // @[RoundAnyRawFNToRecFN.scala 186:16:freechips.rocketchip.system.DefaultRV32Config.fir@173439.4]
  wire [1:0] _T_33; // @[RoundAnyRawFNToRecFN.scala 199:54:freechips.rocketchip.system.DefaultRV32Config.fir@173440.4]
  wire [2:0] _T_34; // @[RoundAnyRawFNToRecFN.scala 199:69:freechips.rocketchip.system.DefaultRV32Config.fir@173441.4]
  wire [9:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@173442.4]
  wire [10:0] sRoundedExp; // @[RoundAnyRawFNToRecFN.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@173442.4]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 202:37:freechips.rocketchip.system.DefaultRV32Config.fir@173443.4]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 206:27:freechips.rocketchip.system.DefaultRV32Config.fir@173446.4]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 256:64:freechips.rocketchip.system.DefaultRV32Config.fir@173474.4]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 259:43:freechips.rocketchip.system.DefaultRV32Config.fir@173478.4]
  wire [8:0] _T_62; // @[RoundAnyRawFNToRecFN.scala 272:18:freechips.rocketchip.system.DefaultRV32Config.fir@173491.4]
  wire [8:0] _T_63; // @[RoundAnyRawFNToRecFN.scala 272:14:freechips.rocketchip.system.DefaultRV32Config.fir@173492.4]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 271:24:freechips.rocketchip.system.DefaultRV32Config.fir@173493.4]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 299:12:freechips.rocketchip.system.DefaultRV32Config.fir@173515.4]
  wire [9:0] _T_88; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@173519.4]
  wire [1:0] _T_90; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@173522.4]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53:freechips.rocketchip.system.DefaultRV32Config.fir@173378.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53:freechips.rocketchip.system.DefaultRV32Config.fir@173380.4]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53:freechips.rocketchip.system.DefaultRV32Config.fir@173381.4]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53:freechips.rocketchip.system.DefaultRV32Config.fir@173382.4]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53:freechips.rocketchip.system.DefaultRV32Config.fir@173383.4]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27:freechips.rocketchip.system.DefaultRV32Config.fir@173384.4]
  assign _T_1 = io_in_sign == 1'h0; // @[RoundAnyRawFNToRecFN.scala 96:66:freechips.rocketchip.system.DefaultRV32Config.fir@173385.4]
  assign _T_2 = roundingMode_max & _T_1; // @[RoundAnyRawFNToRecFN.scala 96:63:freechips.rocketchip.system.DefaultRV32Config.fir@173386.4]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42:freechips.rocketchip.system.DefaultRV32Config.fir@173387.4]
  assign _GEN_0 = {{1{io_in_sExp[7]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@173388.4]
  assign _T_3 = $signed(_GEN_0) + $signed(9'shc0); // @[RoundAnyRawFNToRecFN.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@173388.4]
  assign _T_4 = _T_3[8:0]; // @[RoundAnyRawFNToRecFN.scala 104:14:freechips.rocketchip.system.DefaultRV32Config.fir@173389.4]
  assign sAdjustedExp = {1'b0,$signed(_T_4)}; // @[RoundAnyRawFNToRecFN.scala 104:31:freechips.rocketchip.system.DefaultRV32Config.fir@173390.4]
  assign _T_5 = io_in_sig[32:7]; // @[RoundAnyRawFNToRecFN.scala 115:26:freechips.rocketchip.system.DefaultRV32Config.fir@173391.4]
  assign _T_6 = io_in_sig[6:0]; // @[RoundAnyRawFNToRecFN.scala 116:26:freechips.rocketchip.system.DefaultRV32Config.fir@173392.4]
  assign _T_7 = _T_6 != 7'h0; // @[RoundAnyRawFNToRecFN.scala 116:60:freechips.rocketchip.system.DefaultRV32Config.fir@173393.4]
  assign adjustedSig = {_T_5,_T_7}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@173394.4]
  assign _T_11 = adjustedSig & 27'h2; // @[RoundAnyRawFNToRecFN.scala 173:40:freechips.rocketchip.system.DefaultRV32Config.fir@173413.4]
  assign roundPosBit = _T_11 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 173:56:freechips.rocketchip.system.DefaultRV32Config.fir@173414.4]
  assign _T_12 = adjustedSig & 27'h1; // @[RoundAnyRawFNToRecFN.scala 175:42:freechips.rocketchip.system.DefaultRV32Config.fir@173415.4]
  assign anyRoundExtra = _T_12 != 27'h0; // @[RoundAnyRawFNToRecFN.scala 175:62:freechips.rocketchip.system.DefaultRV32Config.fir@173416.4]
  assign anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 177:36:freechips.rocketchip.system.DefaultRV32Config.fir@173417.4]
  assign _T_13 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 181:38:freechips.rocketchip.system.DefaultRV32Config.fir@173418.4]
  assign _T_14 = _T_13 & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 181:67:freechips.rocketchip.system.DefaultRV32Config.fir@173419.4]
  assign _T_15 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 183:29:freechips.rocketchip.system.DefaultRV32Config.fir@173420.4]
  assign roundIncr = _T_14 | _T_15; // @[RoundAnyRawFNToRecFN.scala 182:31:freechips.rocketchip.system.DefaultRV32Config.fir@173421.4]
  assign _T_16 = adjustedSig | 27'h3; // @[RoundAnyRawFNToRecFN.scala 187:32:freechips.rocketchip.system.DefaultRV32Config.fir@173422.4]
  assign _T_17 = _T_16[26:2]; // @[RoundAnyRawFNToRecFN.scala 187:44:freechips.rocketchip.system.DefaultRV32Config.fir@173423.4]
  assign _T_18 = _T_17 + 25'h1; // @[RoundAnyRawFNToRecFN.scala 187:49:freechips.rocketchip.system.DefaultRV32Config.fir@173424.4]
  assign _T_19 = roundingMode_near_even & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 188:49:freechips.rocketchip.system.DefaultRV32Config.fir@173425.4]
  assign _T_20 = anyRoundExtra == 1'h0; // @[RoundAnyRawFNToRecFN.scala 189:30:freechips.rocketchip.system.DefaultRV32Config.fir@173426.4]
  assign _T_21 = _T_19 & _T_20; // @[RoundAnyRawFNToRecFN.scala 188:64:freechips.rocketchip.system.DefaultRV32Config.fir@173427.4]
  assign _T_23 = _T_21 ? 26'h1 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 188:25:freechips.rocketchip.system.DefaultRV32Config.fir@173429.4]
  assign _T_24 = ~ _T_23; // @[RoundAnyRawFNToRecFN.scala 188:21:freechips.rocketchip.system.DefaultRV32Config.fir@173430.4]
  assign _T_25 = _T_18 & _T_24; // @[RoundAnyRawFNToRecFN.scala 187:61:freechips.rocketchip.system.DefaultRV32Config.fir@173431.4]
  assign _T_27 = adjustedSig & 27'h7fffffc; // @[RoundAnyRawFNToRecFN.scala 193:30:freechips.rocketchip.system.DefaultRV32Config.fir@173433.4]
  assign _T_28 = _T_27[26:2]; // @[RoundAnyRawFNToRecFN.scala 193:43:freechips.rocketchip.system.DefaultRV32Config.fir@173434.4]
  assign _T_29 = roundingMode_odd & anyRound; // @[RoundAnyRawFNToRecFN.scala 194:42:freechips.rocketchip.system.DefaultRV32Config.fir@173435.4]
  assign _T_31 = _T_29 ? 26'h1 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 194:24:freechips.rocketchip.system.DefaultRV32Config.fir@173437.4]
  assign _GEN_1 = {{1'd0}, _T_28}; // @[RoundAnyRawFNToRecFN.scala 193:47:freechips.rocketchip.system.DefaultRV32Config.fir@173438.4]
  assign _T_32 = _GEN_1 | _T_31; // @[RoundAnyRawFNToRecFN.scala 193:47:freechips.rocketchip.system.DefaultRV32Config.fir@173438.4]
  assign roundedSig = roundIncr ? _T_25 : _T_32; // @[RoundAnyRawFNToRecFN.scala 186:16:freechips.rocketchip.system.DefaultRV32Config.fir@173439.4]
  assign _T_33 = roundedSig[25:24]; // @[RoundAnyRawFNToRecFN.scala 199:54:freechips.rocketchip.system.DefaultRV32Config.fir@173440.4]
  assign _T_34 = {1'b0,$signed(_T_33)}; // @[RoundAnyRawFNToRecFN.scala 199:69:freechips.rocketchip.system.DefaultRV32Config.fir@173441.4]
  assign _GEN_2 = {{7{_T_34[2]}},_T_34}; // @[RoundAnyRawFNToRecFN.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@173442.4]
  assign sRoundedExp = $signed(sAdjustedExp) + $signed(_GEN_2); // @[RoundAnyRawFNToRecFN.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@173442.4]
  assign common_expOut = sRoundedExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 202:37:freechips.rocketchip.system.DefaultRV32Config.fir@173443.4]
  assign common_fractOut = roundedSig[22:0]; // @[RoundAnyRawFNToRecFN.scala 206:27:freechips.rocketchip.system.DefaultRV32Config.fir@173446.4]
  assign commonCase = io_in_isZero == 1'h0; // @[RoundAnyRawFNToRecFN.scala 256:64:freechips.rocketchip.system.DefaultRV32Config.fir@173474.4]
  assign inexact = commonCase & anyRound; // @[RoundAnyRawFNToRecFN.scala 259:43:freechips.rocketchip.system.DefaultRV32Config.fir@173478.4]
  assign _T_62 = io_in_isZero ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 272:18:freechips.rocketchip.system.DefaultRV32Config.fir@173491.4]
  assign _T_63 = ~ _T_62; // @[RoundAnyRawFNToRecFN.scala 272:14:freechips.rocketchip.system.DefaultRV32Config.fir@173492.4]
  assign expOut = common_expOut & _T_63; // @[RoundAnyRawFNToRecFN.scala 271:24:freechips.rocketchip.system.DefaultRV32Config.fir@173493.4]
  assign fractOut = io_in_isZero ? 23'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 299:12:freechips.rocketchip.system.DefaultRV32Config.fir@173515.4]
  assign _T_88 = {io_in_sign,expOut}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@173519.4]
  assign _T_90 = {1'h0,inexact}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@173522.4]
  assign io_out = {_T_88,fractOut}; // @[RoundAnyRawFNToRecFN.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@173521.4]
  assign io_exceptionFlags = {3'h0,_T_90}; // @[RoundAnyRawFNToRecFN.scala 306:23:freechips.rocketchip.system.DefaultRV32Config.fir@173526.4]
endmodule

