module DMIToTL( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71022.2]
  input         auto_out_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  output        auto_out_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  output [2:0]  auto_out_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  output [8:0]  auto_out_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  output [3:0]  auto_out_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  output [31:0] auto_out_a_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  output        auto_out_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  input         auto_out_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  input         auto_out_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  input  [31:0] auto_out_d_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  input         auto_out_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71025.4]
  output        io_dmi_req_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
  input         io_dmi_req_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
  input  [6:0]  io_dmi_req_bits_addr, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
  input  [31:0] io_dmi_req_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
  input  [1:0]  io_dmi_req_bits_op, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
  input         io_dmi_resp_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
  output        io_dmi_resp_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
  output [31:0] io_dmi_resp_bits_data, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
  output [1:0]  io_dmi_resp_bits_resp // @[:freechips.rocketchip.system.DefaultRV32Config.fir@71026.4]
);
  wire [8:0] addr; // @[DMI.scala 96:50:freechips.rocketchip.system.DefaultRV32Config.fir@71038.4]
  wire  _T_100; // @[DMI.scala 110:30:freechips.rocketchip.system.DefaultRV32Config.fir@71171.4]
  wire  _T_101; // @[DMI.scala 111:37:freechips.rocketchip.system.DefaultRV32Config.fir@71176.6]
  wire [2:0] _GEN_0; // @[DMI.scala 111:64:freechips.rocketchip.system.DefaultRV32Config.fir@71177.6]
  wire [8:0] _GEN_4; // @[DMI.scala 111:64:freechips.rocketchip.system.DefaultRV32Config.fir@71177.6]
  wire [3:0] _GEN_5; // @[DMI.scala 111:64:freechips.rocketchip.system.DefaultRV32Config.fir@71177.6]
  wire  _T_102; // @[DMI.scala 120:53:freechips.rocketchip.system.DefaultRV32Config.fir@71187.4]
  assign addr = {io_dmi_req_bits_addr, 2'h0}; // @[DMI.scala 96:50:freechips.rocketchip.system.DefaultRV32Config.fir@71038.4]
  assign _T_100 = io_dmi_req_bits_op == 2'h2; // @[DMI.scala 110:30:freechips.rocketchip.system.DefaultRV32Config.fir@71171.4]
  assign _T_101 = io_dmi_req_bits_op == 2'h1; // @[DMI.scala 111:37:freechips.rocketchip.system.DefaultRV32Config.fir@71176.6]
  assign _GEN_0 = _T_101 ? 3'h4 : 3'h1; // @[DMI.scala 111:64:freechips.rocketchip.system.DefaultRV32Config.fir@71177.6]
  assign _GEN_4 = _T_101 ? addr : 9'h40; // @[DMI.scala 111:64:freechips.rocketchip.system.DefaultRV32Config.fir@71177.6]
  assign _GEN_5 = _T_101 ? 4'hf : 4'h0; // @[DMI.scala 111:64:freechips.rocketchip.system.DefaultRV32Config.fir@71177.6]
  assign _T_102 = auto_out_d_bits_corrupt | auto_out_d_bits_denied; // @[DMI.scala 120:53:freechips.rocketchip.system.DefaultRV32Config.fir@71187.4]
  assign auto_out_a_valid = io_dmi_req_valid; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultRV32Config.fir@71034.4]
  assign auto_out_a_bits_opcode = _T_100 ? 3'h0 : _GEN_0; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultRV32Config.fir@71034.4]
  assign auto_out_a_bits_address = _T_100 ? addr : _GEN_4; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultRV32Config.fir@71034.4]
  assign auto_out_a_bits_mask = _T_100 ? 4'hf : _GEN_5; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultRV32Config.fir@71034.4]
  assign auto_out_a_bits_data = _T_100 ? io_dmi_req_bits_data : 32'h0; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultRV32Config.fir@71034.4]
  assign auto_out_d_ready = io_dmi_resp_ready; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultRV32Config.fir@71034.4]
  assign io_dmi_req_ready = auto_out_a_ready; // @[DMI.scala 116:22:freechips.rocketchip.system.DefaultRV32Config.fir@71184.4]
  assign io_dmi_resp_valid = auto_out_d_valid; // @[DMI.scala 118:28:freechips.rocketchip.system.DefaultRV32Config.fir@71185.4]
  assign io_dmi_resp_bits_data = auto_out_d_bits_data; // @[DMI.scala 121:28:freechips.rocketchip.system.DefaultRV32Config.fir@71190.4]
  assign io_dmi_resp_bits_resp = {{1'd0}, _T_102}; // @[DMI.scala 120:28:freechips.rocketchip.system.DefaultRV32Config.fir@71189.4]
endmodule

